magic
tech scmos
timestamp 716090279
<< polycontact >>
rect 0 0 12 4
<< end >>
