magic
tech scmos
timestamp 760840526
<< polysilicon >>
rect 528 56 534 58
rect 528 28 530 56
rect 532 45 534 56
rect 536 56 542 58
rect 536 45 538 56
rect 532 43 538 45
rect 540 45 542 56
rect 544 56 550 58
rect 544 45 546 56
rect 540 43 546 45
rect 548 45 550 56
rect 552 57 558 58
rect 552 53 553 57
rect 557 53 558 57
rect 552 52 558 53
rect 552 48 553 52
rect 557 48 558 52
rect 552 47 558 48
rect 553 45 557 47
rect 548 43 557 45
rect 532 39 538 41
rect 532 28 534 39
rect 528 26 534 28
rect 536 28 538 39
rect 540 39 546 41
rect 540 28 542 39
rect 536 26 542 28
rect 544 28 546 39
rect 548 39 557 41
rect 548 28 550 39
rect 553 37 557 39
rect 544 26 550 28
rect 552 36 558 37
rect 552 32 553 36
rect 557 32 558 36
rect 552 31 558 32
rect 552 27 553 31
rect 557 27 558 31
rect 552 26 558 27
<< metal1 >>
rect 576 81 582 82
rect 576 79 577 81
rect 575 78 577 79
rect 574 77 577 78
rect 581 77 582 81
rect 573 76 582 77
rect 572 75 579 76
rect 571 74 578 75
rect 570 73 577 74
rect 569 72 576 73
rect 568 71 575 72
rect 567 70 574 71
rect 566 69 573 70
rect 565 68 572 69
rect 564 67 571 68
rect 563 66 570 67
rect 562 65 569 66
rect 561 64 568 65
rect 560 63 567 64
rect 559 62 566 63
rect 558 61 565 62
rect 557 60 564 61
rect 556 59 563 60
rect 555 58 562 59
rect 552 57 561 58
rect 552 53 553 57
rect 557 56 560 57
rect 557 55 559 56
rect 557 53 558 55
rect 552 52 558 53
rect 552 48 553 52
rect 557 48 558 52
rect 552 47 558 48
rect 552 36 558 37
rect 552 32 553 36
rect 557 32 558 36
rect 552 31 558 32
rect 552 27 553 31
rect 557 29 558 31
rect 557 28 559 29
rect 557 27 560 28
rect 552 26 561 27
rect 555 25 562 26
rect 556 24 563 25
rect 557 23 564 24
rect 558 22 565 23
rect 559 21 566 22
rect 560 20 567 21
rect 561 19 568 20
rect 562 18 569 19
rect 563 17 570 18
rect 564 16 571 17
rect 565 15 572 16
rect 566 14 573 15
rect 567 13 574 14
rect 568 12 575 13
rect 569 11 576 12
rect 570 10 577 11
rect 571 9 578 10
rect 572 8 579 9
rect 573 7 580 8
rect 574 6 581 7
rect 575 5 582 6
rect 576 4 582 5
rect 577 3 582 4
rect 578 2 582 3
<< metal2 >>
rect 576 81 582 82
rect 576 77 577 81
rect 581 77 582 81
rect 576 76 582 77
<< polycontact >>
rect 553 53 557 57
rect 553 48 557 52
rect 553 32 557 36
rect 553 27 557 31
<< m2contact >>
rect 577 77 581 81
<< substrateopen >>
rect 512 81 572 82
rect 513 80 571 81
rect 514 79 570 80
rect 515 78 569 79
rect 516 77 568 78
rect 517 76 567 77
rect 518 75 566 76
rect 519 74 565 75
rect 520 73 564 74
rect 521 72 563 73
rect 502 71 503 72
rect 522 71 562 72
rect 581 71 582 72
rect 502 70 504 71
rect 523 70 561 71
rect 580 70 582 71
rect 502 69 505 70
rect 524 69 560 70
rect 579 69 582 70
rect 502 68 506 69
rect 525 68 559 69
rect 578 68 582 69
rect 502 67 507 68
rect 526 67 558 68
rect 577 67 582 68
rect 502 66 508 67
rect 527 66 557 67
rect 576 66 582 67
rect 502 65 509 66
rect 528 65 556 66
rect 575 65 582 66
rect 502 64 510 65
rect 529 64 555 65
rect 574 64 582 65
rect 502 63 511 64
rect 530 63 554 64
rect 573 63 582 64
rect 502 62 512 63
rect 572 62 582 63
rect 502 61 513 62
rect 571 61 582 62
rect 502 60 514 61
rect 570 60 582 61
rect 502 59 515 60
rect 569 59 582 60
rect 502 58 516 59
rect 568 58 582 59
rect 502 57 517 58
rect 567 57 582 58
rect 502 56 518 57
rect 566 56 582 57
rect 502 55 519 56
rect 565 55 582 56
rect 502 54 520 55
rect 564 54 582 55
rect 502 30 521 54
rect 563 30 582 54
rect 502 29 520 30
rect 564 29 582 30
rect 502 28 519 29
rect 565 28 582 29
rect 502 27 518 28
rect 566 27 582 28
rect 502 26 517 27
rect 567 26 582 27
rect 502 25 516 26
rect 568 25 582 26
rect 502 24 515 25
rect 569 24 582 25
rect 502 23 514 24
rect 570 23 582 24
rect 502 22 513 23
rect 571 22 582 23
rect 502 21 512 22
rect 572 21 582 22
rect 502 20 511 21
rect 530 20 554 21
rect 573 20 582 21
rect 502 19 510 20
rect 529 19 555 20
rect 574 19 582 20
rect 502 18 509 19
rect 528 18 556 19
rect 575 18 582 19
rect 502 17 508 18
rect 527 17 557 18
rect 576 17 582 18
rect 502 16 507 17
rect 526 16 558 17
rect 577 16 582 17
rect 502 15 506 16
rect 525 15 559 16
rect 578 15 582 16
rect 502 14 505 15
rect 524 14 560 15
rect 579 14 582 15
rect 502 13 504 14
rect 523 13 561 14
rect 580 13 582 14
rect 502 12 503 13
rect 522 12 562 13
rect 581 12 582 13
rect 521 11 563 12
rect 520 10 564 11
rect 519 9 565 10
rect 518 8 566 9
rect 517 7 567 8
rect 516 6 568 7
rect 515 5 569 6
rect 514 4 570 5
rect 513 3 571 4
rect 512 2 572 3
<< pdiffusionstop >>
rect 497 82 587 87
rect 497 2 502 82
rect 582 2 587 82
rect 497 -3 587 2
<< end >>
