magic
tech scmos
timestamp 736072621
<< metal2 >>
rect 1 5 5 16
rect 5 1 6 5
rect 1 0 5 1
<< metal3 >>
rect 0 10 14 16
rect 0 5 14 6
rect 0 1 1 5
rect 5 1 6 5
rect 10 1 14 5
rect 0 0 14 1
<< m3contact >>
rect 1 1 5 5
rect 6 1 10 5
<< end >>
