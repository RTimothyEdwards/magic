magic
tech scmos
timestamp 500617727
<< polysilicon >>
rect -12 6 12 8
<< metal1 >>
rect -12 0 29 3
<< metal2 >>
rect -12 -6 -2 -3
<< labels >>
rlabel polysilicon 11 7 11 7 7 1
rlabel space 11 21 11 21 1 2
rlabel metal1 28 1 28 1 7 5
rlabel space 28 -13 28 -13 5 6
rlabel metal2 -3 -5 -3 -5 7 8
rlabel space 15 -9 15 -9 5 9
rlabel space 5 -21 5 -21 5 10
rlabel space 35 20 35 20 3 3
rlabel space 34 35 34 35 1 4
rlabel space 47 -12 47 -12 3 7
<< end >>
