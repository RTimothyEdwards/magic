magic
tech scmos
timestamp 716915316
<< nwell >>
rect 84 -3742 132 -3710
rect 262 -3741 310 -3698
rect 399 -3741 601 -3698
rect 691 -3741 1070 -3698
rect 1164 -3741 1278 -3698
rect 1362 -3741 1432 -3698
<< metal1 >>
rect -14 -3594 1534 -3586
rect -14 -3846 -6 -3594
rect 0 -3603 80 -3600
rect 0 -3677 3 -3603
rect 77 -3677 80 -3603
rect 114 -3616 125 -3594
rect 118 -3620 121 -3616
rect 114 -3623 125 -3620
rect 118 -3627 121 -3623
rect 114 -3630 125 -3627
rect 118 -3634 121 -3630
rect 160 -3603 240 -3600
rect 0 -3680 80 -3677
rect 76 -3697 80 -3680
rect 160 -3677 163 -3603
rect 237 -3677 240 -3603
rect 160 -3680 240 -3677
rect 320 -3603 400 -3600
rect 320 -3677 323 -3603
rect 397 -3677 400 -3603
rect 434 -3616 445 -3594
rect 438 -3620 441 -3616
rect 434 -3623 445 -3620
rect 438 -3627 441 -3623
rect 434 -3630 445 -3627
rect 438 -3634 441 -3630
rect 480 -3603 560 -3600
rect 320 -3680 400 -3677
rect 480 -3677 483 -3603
rect 557 -3677 560 -3603
rect 480 -3680 560 -3677
rect 640 -3603 720 -3600
rect 640 -3677 643 -3603
rect 717 -3677 720 -3603
rect 754 -3616 765 -3594
rect 758 -3620 761 -3616
rect 754 -3623 765 -3620
rect 758 -3627 761 -3623
rect 754 -3630 765 -3627
rect 758 -3634 761 -3630
rect 800 -3603 880 -3600
rect 640 -3680 720 -3677
rect 800 -3677 803 -3603
rect 877 -3677 880 -3603
rect 800 -3680 880 -3677
rect 960 -3603 1040 -3600
rect 960 -3677 963 -3603
rect 1037 -3675 1040 -3603
rect 1074 -3616 1085 -3594
rect 1078 -3620 1081 -3616
rect 1074 -3623 1085 -3620
rect 1078 -3627 1081 -3623
rect 1074 -3630 1085 -3627
rect 1078 -3634 1081 -3630
rect 1120 -3603 1200 -3600
rect 1037 -3677 1060 -3675
rect 960 -3680 1060 -3677
rect 1120 -3677 1123 -3603
rect 1197 -3677 1200 -3603
rect 1120 -3680 1200 -3677
rect 1280 -3603 1360 -3600
rect 1280 -3677 1283 -3603
rect 1357 -3677 1360 -3603
rect 1394 -3616 1405 -3594
rect 1475 -3600 1486 -3594
rect 1398 -3620 1401 -3616
rect 1394 -3623 1405 -3620
rect 1398 -3627 1401 -3623
rect 1394 -3630 1405 -3627
rect 1398 -3634 1401 -3630
rect 1440 -3603 1520 -3600
rect 1280 -3680 1360 -3677
rect 1440 -3677 1443 -3603
rect 1517 -3677 1520 -3603
rect 1440 -3680 1520 -3677
rect 160 -3697 164 -3680
rect 320 -3682 325 -3680
rect 76 -3701 112 -3697
rect 85 -3716 89 -3715
rect 108 -3718 112 -3701
rect 106 -3724 112 -3718
rect 110 -3728 112 -3724
rect 115 -3701 164 -3697
rect 288 -3687 325 -3682
rect 263 -3700 269 -3699
rect 115 -3721 119 -3701
rect 127 -3716 131 -3715
rect 115 -3724 121 -3721
rect 115 -3728 117 -3724
rect 95 -3731 99 -3728
rect 115 -3731 121 -3728
rect 95 -3734 121 -3731
rect 85 -3737 89 -3736
rect 127 -3737 131 -3736
rect 85 -3741 86 -3737
rect 130 -3741 164 -3737
rect 267 -3703 269 -3700
rect 288 -3708 292 -3687
rect 480 -3690 485 -3680
rect 640 -3687 645 -3680
rect 284 -3712 292 -3708
rect 295 -3695 485 -3690
rect 596 -3692 645 -3687
rect 872 -3686 880 -3680
rect 273 -3714 277 -3712
rect 273 -3730 277 -3726
rect 284 -3723 288 -3716
rect 295 -3714 299 -3695
rect 596 -3699 600 -3692
rect 872 -3693 1052 -3686
rect 302 -3703 303 -3699
rect 307 -3703 309 -3699
rect 295 -3730 299 -3726
rect 273 -3733 299 -3730
rect 305 -3706 309 -3703
rect 305 -3736 309 -3734
rect 267 -3740 268 -3736
rect 308 -3740 309 -3736
rect 400 -3700 406 -3699
rect 404 -3703 406 -3700
rect 594 -3703 596 -3699
rect 410 -3709 590 -3706
rect 410 -3714 414 -3709
rect 410 -3727 414 -3726
rect 421 -3723 425 -3716
rect 432 -3714 436 -3709
rect 432 -3727 436 -3726
rect 443 -3723 447 -3716
rect 454 -3714 458 -3709
rect 454 -3727 458 -3726
rect 465 -3723 469 -3716
rect 476 -3714 480 -3709
rect 476 -3727 480 -3726
rect 487 -3723 491 -3716
rect 498 -3714 502 -3709
rect 498 -3727 502 -3726
rect 509 -3723 513 -3716
rect 520 -3714 524 -3709
rect 520 -3727 524 -3726
rect 531 -3723 535 -3716
rect 542 -3714 546 -3709
rect 542 -3727 546 -3726
rect 553 -3723 557 -3716
rect 564 -3714 568 -3709
rect 564 -3727 568 -3726
rect 575 -3723 579 -3716
rect 421 -3730 425 -3727
rect 443 -3730 447 -3727
rect 465 -3730 469 -3727
rect 487 -3730 491 -3727
rect 509 -3730 513 -3727
rect 531 -3730 535 -3727
rect 553 -3730 557 -3727
rect 575 -3730 579 -3727
rect 586 -3714 590 -3709
rect 421 -3733 583 -3730
rect 404 -3740 406 -3736
rect 574 -3740 575 -3736
rect 160 -3760 164 -3741
rect 305 -3748 309 -3740
rect 305 -3753 400 -3748
rect 395 -3760 400 -3753
rect 579 -3755 583 -3733
rect 556 -3760 583 -3755
rect 586 -3755 590 -3726
rect 596 -3736 600 -3735
rect 593 -3740 594 -3736
rect 598 -3740 600 -3736
rect 692 -3700 697 -3699
rect 696 -3703 697 -3700
rect 1048 -3706 1052 -3693
rect 713 -3709 1052 -3706
rect 713 -3712 717 -3709
rect 735 -3712 739 -3709
rect 757 -3712 761 -3709
rect 779 -3712 783 -3709
rect 801 -3712 805 -3709
rect 823 -3712 827 -3709
rect 845 -3712 849 -3709
rect 867 -3712 871 -3709
rect 889 -3712 893 -3709
rect 911 -3712 915 -3709
rect 933 -3712 937 -3709
rect 955 -3712 959 -3709
rect 978 -3712 982 -3709
rect 1000 -3712 1004 -3709
rect 1022 -3712 1026 -3709
rect 1044 -3712 1048 -3709
rect 702 -3714 706 -3712
rect 702 -3730 706 -3726
rect 713 -3723 717 -3716
rect 724 -3714 728 -3712
rect 724 -3730 728 -3726
rect 735 -3723 739 -3716
rect 746 -3714 750 -3712
rect 746 -3730 750 -3726
rect 757 -3723 761 -3716
rect 768 -3714 772 -3712
rect 768 -3730 772 -3726
rect 779 -3723 783 -3716
rect 790 -3714 794 -3712
rect 790 -3730 794 -3726
rect 801 -3723 805 -3716
rect 812 -3714 816 -3712
rect 812 -3730 816 -3726
rect 823 -3723 827 -3716
rect 834 -3714 838 -3712
rect 834 -3730 838 -3726
rect 845 -3723 849 -3716
rect 856 -3714 860 -3712
rect 856 -3730 860 -3726
rect 867 -3723 871 -3716
rect 878 -3714 882 -3712
rect 878 -3730 882 -3726
rect 889 -3723 893 -3716
rect 900 -3714 904 -3712
rect 900 -3730 904 -3726
rect 911 -3723 915 -3716
rect 922 -3714 926 -3712
rect 922 -3730 926 -3726
rect 933 -3723 937 -3716
rect 944 -3714 948 -3712
rect 944 -3730 948 -3726
rect 955 -3723 959 -3716
rect 966 -3714 970 -3712
rect 966 -3730 970 -3726
rect 978 -3723 982 -3716
rect 989 -3714 993 -3712
rect 989 -3730 993 -3726
rect 1000 -3723 1004 -3716
rect 1011 -3714 1015 -3712
rect 1011 -3730 1015 -3726
rect 1022 -3723 1026 -3716
rect 1033 -3714 1037 -3712
rect 1033 -3730 1037 -3726
rect 1044 -3723 1048 -3716
rect 1055 -3714 1060 -3680
rect 1195 -3699 1200 -3680
rect 1355 -3699 1360 -3680
rect 1063 -3703 1064 -3699
rect 1068 -3703 1069 -3699
rect 1059 -3726 1060 -3714
rect 1055 -3730 1060 -3726
rect 702 -3733 1060 -3730
rect 1065 -3704 1069 -3703
rect 696 -3740 698 -3736
rect 1062 -3740 1065 -3736
rect 1169 -3703 1171 -3699
rect 1275 -3703 1277 -3699
rect 1273 -3706 1277 -3703
rect 1355 -3700 1369 -3699
rect 1355 -3705 1363 -3700
rect 1165 -3736 1169 -3735
rect 1175 -3709 1267 -3706
rect 1175 -3714 1179 -3709
rect 1165 -3740 1166 -3736
rect 1170 -3740 1172 -3736
rect 586 -3760 644 -3755
rect 872 -3760 880 -3740
rect 1175 -3749 1179 -3726
rect 1186 -3723 1190 -3716
rect 1197 -3714 1201 -3709
rect 1197 -3727 1201 -3726
rect 1208 -3723 1212 -3716
rect 1219 -3714 1223 -3709
rect 1219 -3727 1223 -3726
rect 1230 -3723 1234 -3716
rect 1241 -3714 1245 -3709
rect 1241 -3727 1245 -3726
rect 1252 -3723 1256 -3716
rect 1263 -3714 1267 -3709
rect 1263 -3727 1267 -3726
rect 1186 -3730 1190 -3727
rect 1208 -3730 1212 -3727
rect 1230 -3730 1234 -3727
rect 1252 -3730 1256 -3727
rect 1035 -3754 1179 -3749
rect 1182 -3733 1256 -3730
rect 1035 -3760 1040 -3754
rect 1182 -3760 1186 -3733
rect 1273 -3736 1277 -3734
rect 1367 -3703 1369 -3700
rect 1425 -3703 1427 -3699
rect 1373 -3709 1421 -3706
rect 1373 -3714 1377 -3709
rect 1373 -3727 1377 -3726
rect 1384 -3723 1388 -3716
rect 1395 -3714 1399 -3709
rect 1395 -3727 1399 -3726
rect 1406 -3723 1410 -3716
rect 1384 -3730 1388 -3727
rect 1406 -3730 1410 -3727
rect 1417 -3714 1421 -3709
rect 1384 -3733 1414 -3730
rect 1367 -3740 1369 -3736
rect 1405 -3740 1407 -3736
rect 1410 -3749 1414 -3733
rect 1355 -3753 1414 -3749
rect 1417 -3749 1421 -3726
rect 1427 -3736 1431 -3735
rect 1424 -3740 1425 -3736
rect 1429 -3740 1431 -3736
rect 1417 -3753 1445 -3749
rect 1355 -3760 1360 -3753
rect 0 -3763 80 -3760
rect 0 -3837 3 -3763
rect 77 -3837 80 -3763
rect 0 -3840 80 -3837
rect 160 -3763 240 -3760
rect 160 -3837 163 -3763
rect 237 -3837 240 -3763
rect 320 -3763 400 -3760
rect 160 -3840 240 -3837
rect 278 -3810 281 -3806
rect 274 -3813 285 -3810
rect 278 -3817 281 -3813
rect 274 -3820 285 -3817
rect 278 -3824 281 -3820
rect 35 -3846 46 -3840
rect 274 -3846 285 -3824
rect 320 -3837 323 -3763
rect 397 -3837 400 -3763
rect 320 -3840 400 -3837
rect 480 -3763 560 -3760
rect 480 -3837 483 -3763
rect 557 -3837 560 -3763
rect 640 -3763 720 -3760
rect 480 -3840 560 -3837
rect 598 -3810 601 -3806
rect 594 -3813 605 -3810
rect 598 -3817 601 -3813
rect 594 -3820 605 -3817
rect 598 -3824 601 -3820
rect 594 -3846 605 -3824
rect 640 -3837 643 -3763
rect 717 -3837 720 -3763
rect 640 -3840 720 -3837
rect 800 -3763 880 -3760
rect 800 -3837 803 -3763
rect 877 -3837 880 -3763
rect 960 -3763 1040 -3760
rect 800 -3840 880 -3837
rect 918 -3810 921 -3806
rect 914 -3813 925 -3810
rect 918 -3817 921 -3813
rect 914 -3820 925 -3817
rect 918 -3824 921 -3820
rect 914 -3846 925 -3824
rect 960 -3837 963 -3763
rect 1037 -3837 1040 -3763
rect 960 -3840 1040 -3837
rect 1120 -3763 1200 -3760
rect 1120 -3837 1123 -3763
rect 1197 -3837 1200 -3763
rect 1280 -3763 1360 -3760
rect 1120 -3840 1200 -3837
rect 1238 -3810 1241 -3806
rect 1234 -3813 1245 -3810
rect 1238 -3817 1241 -3813
rect 1234 -3820 1245 -3817
rect 1238 -3824 1241 -3820
rect 1234 -3846 1245 -3824
rect 1280 -3837 1283 -3763
rect 1357 -3837 1360 -3763
rect 1280 -3840 1360 -3837
rect 1440 -3760 1445 -3753
rect 1440 -3763 1520 -3760
rect 1440 -3837 1443 -3763
rect 1517 -3837 1520 -3763
rect 1440 -3840 1520 -3837
rect 1526 -3846 1534 -3594
rect -14 -3854 1534 -3846
<< metal2 >>
rect 0 -3603 80 -3600
rect 0 -3677 3 -3603
rect 77 -3677 80 -3603
rect 0 -3680 80 -3677
rect 160 -3603 240 -3600
rect 160 -3677 163 -3603
rect 237 -3677 240 -3603
rect 160 -3680 240 -3677
rect 320 -3603 400 -3600
rect 320 -3677 323 -3603
rect 397 -3677 400 -3603
rect 320 -3680 400 -3677
rect 480 -3603 560 -3600
rect 480 -3677 483 -3603
rect 557 -3677 560 -3603
rect 480 -3680 560 -3677
rect 640 -3603 720 -3600
rect 640 -3677 643 -3603
rect 717 -3677 720 -3603
rect 640 -3680 720 -3677
rect 800 -3603 880 -3600
rect 800 -3677 803 -3603
rect 877 -3677 880 -3603
rect 800 -3680 880 -3677
rect 960 -3603 1040 -3600
rect 960 -3677 963 -3603
rect 1037 -3677 1040 -3603
rect 960 -3680 1040 -3677
rect 1120 -3603 1200 -3600
rect 1120 -3677 1123 -3603
rect 1197 -3677 1200 -3603
rect 1120 -3680 1200 -3677
rect 1280 -3603 1360 -3600
rect 1280 -3677 1283 -3603
rect 1357 -3677 1360 -3603
rect 1280 -3680 1360 -3677
rect 1440 -3603 1520 -3600
rect 1440 -3677 1443 -3603
rect 1517 -3677 1520 -3603
rect 1440 -3680 1520 -3677
rect 0 -3763 80 -3760
rect 0 -3837 3 -3763
rect 77 -3837 80 -3763
rect 0 -3840 80 -3837
rect 160 -3763 240 -3760
rect 160 -3837 163 -3763
rect 237 -3837 240 -3763
rect 160 -3840 240 -3837
rect 320 -3763 400 -3760
rect 320 -3837 323 -3763
rect 397 -3837 400 -3763
rect 320 -3840 400 -3837
rect 480 -3763 560 -3760
rect 480 -3837 483 -3763
rect 557 -3837 560 -3763
rect 480 -3840 560 -3837
rect 640 -3763 720 -3760
rect 640 -3837 643 -3763
rect 717 -3837 720 -3763
rect 640 -3840 720 -3837
rect 800 -3763 880 -3760
rect 800 -3837 803 -3763
rect 877 -3837 880 -3763
rect 800 -3840 880 -3837
rect 960 -3763 1040 -3760
rect 960 -3837 963 -3763
rect 1037 -3837 1040 -3763
rect 960 -3840 1040 -3837
rect 1120 -3763 1200 -3760
rect 1120 -3837 1123 -3763
rect 1197 -3837 1200 -3763
rect 1120 -3840 1200 -3837
rect 1280 -3763 1360 -3760
rect 1280 -3837 1283 -3763
rect 1357 -3837 1360 -3763
rect 1280 -3840 1360 -3837
rect 1440 -3763 1520 -3760
rect 1440 -3837 1443 -3763
rect 1517 -3837 1520 -3763
rect 1440 -3840 1520 -3837
<< collector >>
rect 262 -3699 310 -3698
rect 262 -3700 269 -3699
rect 84 -3711 132 -3710
rect 84 -3715 85 -3711
rect 105 -3715 122 -3711
rect 131 -3715 132 -3711
rect 84 -3716 132 -3715
rect 84 -3736 85 -3716
rect 89 -3736 90 -3716
rect 126 -3736 127 -3716
rect 131 -3736 132 -3716
rect 84 -3737 132 -3736
rect 84 -3741 86 -3737
rect 130 -3741 132 -3737
rect 262 -3740 263 -3700
rect 267 -3703 269 -3700
rect 285 -3703 303 -3699
rect 307 -3703 310 -3699
rect 267 -3704 310 -3703
rect 267 -3735 268 -3704
rect 304 -3706 310 -3704
rect 304 -3734 305 -3706
rect 309 -3734 310 -3706
rect 304 -3735 310 -3734
rect 267 -3736 310 -3735
rect 267 -3740 268 -3736
rect 308 -3740 310 -3736
rect 262 -3741 310 -3740
rect 399 -3699 601 -3698
rect 399 -3700 406 -3699
rect 399 -3740 400 -3700
rect 404 -3703 406 -3700
rect 594 -3703 596 -3699
rect 404 -3704 596 -3703
rect 404 -3735 405 -3704
rect 595 -3735 596 -3704
rect 600 -3735 601 -3699
rect 404 -3736 601 -3735
rect 404 -3740 406 -3736
rect 574 -3740 594 -3736
rect 598 -3740 601 -3736
rect 399 -3741 601 -3740
rect 691 -3699 1070 -3698
rect 691 -3700 697 -3699
rect 691 -3740 692 -3700
rect 696 -3703 697 -3700
rect 1045 -3703 1064 -3699
rect 1068 -3703 1070 -3699
rect 696 -3704 1070 -3703
rect 696 -3735 697 -3704
rect 1064 -3735 1065 -3704
rect 696 -3736 1065 -3735
rect 696 -3740 698 -3736
rect 1062 -3740 1065 -3736
rect 1069 -3740 1070 -3704
rect 691 -3741 1070 -3740
rect 1164 -3699 1278 -3698
rect 1164 -3735 1165 -3699
rect 1169 -3703 1171 -3699
rect 1275 -3703 1278 -3699
rect 1169 -3704 1278 -3703
rect 1169 -3735 1170 -3704
rect 1272 -3706 1278 -3704
rect 1272 -3734 1273 -3706
rect 1277 -3734 1278 -3706
rect 1272 -3735 1278 -3734
rect 1164 -3736 1278 -3735
rect 1164 -3740 1166 -3736
rect 1170 -3740 1189 -3736
rect 1277 -3740 1278 -3736
rect 1164 -3741 1278 -3740
rect 1362 -3699 1432 -3698
rect 1362 -3700 1369 -3699
rect 1362 -3740 1363 -3700
rect 1367 -3703 1369 -3700
rect 1425 -3703 1427 -3699
rect 1367 -3704 1427 -3703
rect 1367 -3735 1368 -3704
rect 1426 -3735 1427 -3704
rect 1431 -3735 1432 -3699
rect 1367 -3736 1432 -3735
rect 1367 -3740 1369 -3736
rect 1405 -3740 1425 -3736
rect 1429 -3740 1432 -3736
rect 1362 -3741 1432 -3740
rect 84 -3742 132 -3741
<< pbase >>
rect 94 -3724 122 -3720
rect 94 -3728 95 -3724
rect 99 -3728 106 -3724
rect 110 -3728 117 -3724
rect 121 -3728 122 -3724
rect 94 -3732 122 -3728
rect 272 -3712 300 -3708
rect 272 -3714 284 -3712
rect 272 -3726 273 -3714
rect 277 -3716 284 -3714
rect 288 -3714 300 -3712
rect 288 -3716 295 -3714
rect 277 -3723 295 -3716
rect 277 -3726 284 -3723
rect 272 -3727 284 -3726
rect 288 -3726 295 -3723
rect 299 -3726 300 -3714
rect 288 -3727 300 -3726
rect 272 -3731 300 -3727
rect 409 -3712 591 -3708
rect 409 -3714 421 -3712
rect 409 -3726 410 -3714
rect 414 -3716 421 -3714
rect 425 -3714 443 -3712
rect 425 -3716 432 -3714
rect 414 -3723 432 -3716
rect 414 -3726 421 -3723
rect 409 -3727 421 -3726
rect 425 -3726 432 -3723
rect 436 -3716 443 -3714
rect 447 -3714 465 -3712
rect 447 -3716 454 -3714
rect 436 -3723 454 -3716
rect 436 -3726 443 -3723
rect 425 -3727 443 -3726
rect 447 -3726 454 -3723
rect 458 -3716 465 -3714
rect 469 -3714 487 -3712
rect 469 -3716 476 -3714
rect 458 -3723 476 -3716
rect 458 -3726 465 -3723
rect 447 -3727 465 -3726
rect 469 -3726 476 -3723
rect 480 -3716 487 -3714
rect 491 -3714 509 -3712
rect 491 -3716 498 -3714
rect 480 -3723 498 -3716
rect 480 -3726 487 -3723
rect 469 -3727 487 -3726
rect 491 -3726 498 -3723
rect 502 -3716 509 -3714
rect 513 -3714 531 -3712
rect 513 -3716 520 -3714
rect 502 -3723 520 -3716
rect 502 -3726 509 -3723
rect 491 -3727 509 -3726
rect 513 -3726 520 -3723
rect 524 -3716 531 -3714
rect 535 -3714 553 -3712
rect 535 -3716 542 -3714
rect 524 -3723 542 -3716
rect 524 -3726 531 -3723
rect 513 -3727 531 -3726
rect 535 -3726 542 -3723
rect 546 -3716 553 -3714
rect 557 -3714 575 -3712
rect 557 -3716 564 -3714
rect 546 -3723 564 -3716
rect 546 -3726 553 -3723
rect 535 -3727 553 -3726
rect 557 -3726 564 -3723
rect 568 -3716 575 -3714
rect 579 -3714 591 -3712
rect 579 -3716 586 -3714
rect 568 -3723 586 -3716
rect 568 -3726 575 -3723
rect 557 -3727 575 -3726
rect 579 -3726 586 -3723
rect 590 -3726 591 -3714
rect 579 -3727 591 -3726
rect 409 -3731 591 -3727
rect 701 -3712 1060 -3708
rect 701 -3714 713 -3712
rect 701 -3726 702 -3714
rect 706 -3716 713 -3714
rect 717 -3714 735 -3712
rect 717 -3716 724 -3714
rect 706 -3723 724 -3716
rect 706 -3726 713 -3723
rect 701 -3727 713 -3726
rect 717 -3726 724 -3723
rect 728 -3716 735 -3714
rect 739 -3714 757 -3712
rect 739 -3716 746 -3714
rect 728 -3723 746 -3716
rect 728 -3726 735 -3723
rect 717 -3727 735 -3726
rect 739 -3726 746 -3723
rect 750 -3716 757 -3714
rect 761 -3714 779 -3712
rect 761 -3716 768 -3714
rect 750 -3723 768 -3716
rect 750 -3726 757 -3723
rect 739 -3727 757 -3726
rect 761 -3726 768 -3723
rect 772 -3716 779 -3714
rect 783 -3714 801 -3712
rect 783 -3716 790 -3714
rect 772 -3723 790 -3716
rect 772 -3726 779 -3723
rect 761 -3727 779 -3726
rect 783 -3726 790 -3723
rect 794 -3716 801 -3714
rect 805 -3714 823 -3712
rect 805 -3716 812 -3714
rect 794 -3723 812 -3716
rect 794 -3726 801 -3723
rect 783 -3727 801 -3726
rect 805 -3726 812 -3723
rect 816 -3716 823 -3714
rect 827 -3714 845 -3712
rect 827 -3716 834 -3714
rect 816 -3723 834 -3716
rect 816 -3726 823 -3723
rect 805 -3727 823 -3726
rect 827 -3726 834 -3723
rect 838 -3716 845 -3714
rect 849 -3714 867 -3712
rect 849 -3716 856 -3714
rect 838 -3723 856 -3716
rect 838 -3726 845 -3723
rect 827 -3727 845 -3726
rect 849 -3726 856 -3723
rect 860 -3716 867 -3714
rect 871 -3714 889 -3712
rect 871 -3716 878 -3714
rect 860 -3723 878 -3716
rect 860 -3726 867 -3723
rect 849 -3727 867 -3726
rect 871 -3726 878 -3723
rect 882 -3716 889 -3714
rect 893 -3714 911 -3712
rect 893 -3716 900 -3714
rect 882 -3723 900 -3716
rect 882 -3726 889 -3723
rect 871 -3727 889 -3726
rect 893 -3726 900 -3723
rect 904 -3716 911 -3714
rect 915 -3714 933 -3712
rect 915 -3716 922 -3714
rect 904 -3723 922 -3716
rect 904 -3726 911 -3723
rect 893 -3727 911 -3726
rect 915 -3726 922 -3723
rect 926 -3716 933 -3714
rect 937 -3714 955 -3712
rect 937 -3716 944 -3714
rect 926 -3723 944 -3716
rect 926 -3726 933 -3723
rect 915 -3727 933 -3726
rect 937 -3726 944 -3723
rect 948 -3716 955 -3714
rect 959 -3714 978 -3712
rect 959 -3716 966 -3714
rect 948 -3723 966 -3716
rect 948 -3726 955 -3723
rect 937 -3727 955 -3726
rect 959 -3726 966 -3723
rect 970 -3716 978 -3714
rect 982 -3714 1000 -3712
rect 982 -3716 989 -3714
rect 970 -3723 989 -3716
rect 970 -3726 978 -3723
rect 959 -3727 978 -3726
rect 982 -3726 989 -3723
rect 993 -3716 1000 -3714
rect 1004 -3714 1022 -3712
rect 1004 -3716 1011 -3714
rect 993 -3723 1011 -3716
rect 993 -3726 1000 -3723
rect 982 -3727 1000 -3726
rect 1004 -3726 1011 -3723
rect 1015 -3716 1022 -3714
rect 1026 -3714 1044 -3712
rect 1026 -3716 1033 -3714
rect 1015 -3723 1033 -3716
rect 1015 -3726 1022 -3723
rect 1004 -3727 1022 -3726
rect 1026 -3726 1033 -3723
rect 1037 -3716 1044 -3714
rect 1048 -3714 1060 -3712
rect 1048 -3716 1055 -3714
rect 1037 -3723 1055 -3716
rect 1037 -3726 1044 -3723
rect 1026 -3727 1044 -3726
rect 1048 -3726 1055 -3723
rect 1059 -3726 1060 -3714
rect 1048 -3727 1060 -3726
rect 701 -3731 1060 -3727
rect 1174 -3712 1268 -3708
rect 1174 -3714 1186 -3712
rect 1174 -3726 1175 -3714
rect 1179 -3716 1186 -3714
rect 1190 -3714 1208 -3712
rect 1190 -3716 1197 -3714
rect 1179 -3723 1197 -3716
rect 1179 -3726 1186 -3723
rect 1174 -3727 1186 -3726
rect 1190 -3726 1197 -3723
rect 1201 -3716 1208 -3714
rect 1212 -3714 1230 -3712
rect 1212 -3716 1219 -3714
rect 1201 -3723 1219 -3716
rect 1201 -3726 1208 -3723
rect 1190 -3727 1208 -3726
rect 1212 -3726 1219 -3723
rect 1223 -3716 1230 -3714
rect 1234 -3714 1252 -3712
rect 1234 -3716 1241 -3714
rect 1223 -3723 1241 -3716
rect 1223 -3726 1230 -3723
rect 1212 -3727 1230 -3726
rect 1234 -3726 1241 -3723
rect 1245 -3716 1252 -3714
rect 1256 -3714 1268 -3712
rect 1256 -3716 1263 -3714
rect 1245 -3723 1263 -3716
rect 1245 -3726 1252 -3723
rect 1234 -3727 1252 -3726
rect 1256 -3726 1263 -3723
rect 1267 -3726 1268 -3714
rect 1256 -3727 1268 -3726
rect 1174 -3731 1268 -3727
rect 1372 -3712 1422 -3708
rect 1372 -3714 1384 -3712
rect 1372 -3726 1373 -3714
rect 1377 -3716 1384 -3714
rect 1388 -3714 1406 -3712
rect 1388 -3716 1395 -3714
rect 1377 -3723 1395 -3716
rect 1377 -3726 1384 -3723
rect 1372 -3727 1384 -3726
rect 1388 -3726 1395 -3723
rect 1399 -3716 1406 -3714
rect 1410 -3714 1422 -3712
rect 1410 -3716 1417 -3714
rect 1399 -3723 1417 -3716
rect 1399 -3726 1406 -3723
rect 1388 -3727 1406 -3726
rect 1410 -3726 1417 -3723
rect 1421 -3726 1422 -3714
rect 1410 -3727 1422 -3726
rect 1372 -3731 1422 -3727
<< collectorcontact >>
rect 85 -3715 105 -3711
rect 122 -3715 131 -3711
rect 85 -3736 89 -3716
rect 127 -3736 131 -3716
rect 86 -3741 130 -3737
rect 263 -3740 267 -3700
rect 269 -3703 285 -3699
rect 303 -3703 307 -3699
rect 305 -3734 309 -3706
rect 268 -3740 308 -3736
rect 400 -3740 404 -3700
rect 406 -3703 594 -3699
rect 596 -3735 600 -3699
rect 406 -3740 574 -3736
rect 594 -3740 598 -3736
rect 692 -3740 696 -3700
rect 697 -3703 1045 -3699
rect 1064 -3703 1068 -3699
rect 698 -3740 1062 -3736
rect 1065 -3740 1069 -3704
rect 1165 -3735 1169 -3699
rect 1171 -3703 1275 -3699
rect 1273 -3734 1277 -3706
rect 1166 -3740 1170 -3736
rect 1189 -3740 1277 -3736
rect 1363 -3740 1367 -3700
rect 1369 -3703 1425 -3699
rect 1427 -3735 1431 -3699
rect 1369 -3740 1405 -3736
rect 1425 -3740 1429 -3736
<< emittercontact >>
rect 106 -3728 110 -3724
rect 284 -3716 288 -3712
rect 284 -3727 288 -3723
rect 421 -3716 425 -3712
rect 421 -3727 425 -3723
rect 443 -3716 447 -3712
rect 443 -3727 447 -3723
rect 465 -3716 469 -3712
rect 465 -3727 469 -3723
rect 487 -3716 491 -3712
rect 487 -3727 491 -3723
rect 509 -3716 513 -3712
rect 509 -3727 513 -3723
rect 531 -3716 535 -3712
rect 531 -3727 535 -3723
rect 553 -3716 557 -3712
rect 553 -3727 557 -3723
rect 575 -3716 579 -3712
rect 575 -3727 579 -3723
rect 713 -3716 717 -3712
rect 713 -3727 717 -3723
rect 735 -3716 739 -3712
rect 735 -3727 739 -3723
rect 757 -3716 761 -3712
rect 757 -3727 761 -3723
rect 779 -3716 783 -3712
rect 779 -3727 783 -3723
rect 801 -3716 805 -3712
rect 801 -3727 805 -3723
rect 823 -3716 827 -3712
rect 823 -3727 827 -3723
rect 845 -3716 849 -3712
rect 845 -3727 849 -3723
rect 867 -3716 871 -3712
rect 867 -3727 871 -3723
rect 889 -3716 893 -3712
rect 889 -3727 893 -3723
rect 911 -3716 915 -3712
rect 911 -3727 915 -3723
rect 933 -3716 937 -3712
rect 933 -3727 937 -3723
rect 955 -3716 959 -3712
rect 955 -3727 959 -3723
rect 978 -3716 982 -3712
rect 978 -3727 982 -3723
rect 1000 -3716 1004 -3712
rect 1000 -3727 1004 -3723
rect 1022 -3716 1026 -3712
rect 1022 -3727 1026 -3723
rect 1044 -3716 1048 -3712
rect 1044 -3727 1048 -3723
rect 1186 -3716 1190 -3712
rect 1186 -3727 1190 -3723
rect 1208 -3716 1212 -3712
rect 1208 -3727 1212 -3723
rect 1230 -3716 1234 -3712
rect 1230 -3727 1234 -3723
rect 1252 -3716 1256 -3712
rect 1252 -3727 1256 -3723
rect 1384 -3716 1388 -3712
rect 1384 -3727 1388 -3723
rect 1406 -3716 1410 -3712
rect 1406 -3727 1410 -3723
<< pbasecontact >>
rect 95 -3728 99 -3724
rect 117 -3728 121 -3724
rect 273 -3726 277 -3714
rect 295 -3726 299 -3714
rect 410 -3726 414 -3714
rect 432 -3726 436 -3714
rect 454 -3726 458 -3714
rect 476 -3726 480 -3714
rect 498 -3726 502 -3714
rect 520 -3726 524 -3714
rect 542 -3726 546 -3714
rect 564 -3726 568 -3714
rect 586 -3726 590 -3714
rect 702 -3726 706 -3714
rect 724 -3726 728 -3714
rect 746 -3726 750 -3714
rect 768 -3726 772 -3714
rect 790 -3726 794 -3714
rect 812 -3726 816 -3714
rect 834 -3726 838 -3714
rect 856 -3726 860 -3714
rect 878 -3726 882 -3714
rect 900 -3726 904 -3714
rect 922 -3726 926 -3714
rect 944 -3726 948 -3714
rect 966 -3726 970 -3714
rect 989 -3726 993 -3714
rect 1011 -3726 1015 -3714
rect 1033 -3726 1037 -3714
rect 1055 -3726 1059 -3714
rect 1175 -3726 1179 -3714
rect 1197 -3726 1201 -3714
rect 1219 -3726 1223 -3714
rect 1241 -3726 1245 -3714
rect 1263 -3726 1267 -3714
rect 1373 -3726 1377 -3714
rect 1395 -3726 1399 -3714
rect 1417 -3726 1421 -3714
<< m2contact >>
rect 3 -3677 77 -3603
rect 163 -3677 237 -3603
rect 323 -3677 397 -3603
rect 483 -3677 557 -3603
rect 643 -3677 717 -3603
rect 803 -3677 877 -3603
rect 963 -3677 1037 -3603
rect 1123 -3677 1197 -3603
rect 1283 -3677 1357 -3603
rect 1443 -3677 1517 -3603
rect 3 -3837 77 -3763
rect 163 -3837 237 -3763
rect 323 -3837 397 -3763
rect 483 -3837 557 -3763
rect 643 -3837 717 -3763
rect 803 -3837 877 -3763
rect 963 -3837 1037 -3763
rect 1123 -3837 1197 -3763
rect 1283 -3837 1357 -3763
rect 1443 -3837 1517 -3763
<< psubstratepcontact >>
rect 114 -3620 118 -3616
rect 121 -3620 125 -3616
rect 114 -3627 118 -3623
rect 121 -3627 125 -3623
rect 114 -3634 118 -3630
rect 121 -3634 125 -3630
rect 434 -3620 438 -3616
rect 441 -3620 445 -3616
rect 434 -3627 438 -3623
rect 441 -3627 445 -3623
rect 434 -3634 438 -3630
rect 441 -3634 445 -3630
rect 754 -3620 758 -3616
rect 761 -3620 765 -3616
rect 754 -3627 758 -3623
rect 761 -3627 765 -3623
rect 754 -3634 758 -3630
rect 761 -3634 765 -3630
rect 1074 -3620 1078 -3616
rect 1081 -3620 1085 -3616
rect 1074 -3627 1078 -3623
rect 1081 -3627 1085 -3623
rect 1074 -3634 1078 -3630
rect 1081 -3634 1085 -3630
rect 1394 -3620 1398 -3616
rect 1401 -3620 1405 -3616
rect 1394 -3627 1398 -3623
rect 1401 -3627 1405 -3623
rect 1394 -3634 1398 -3630
rect 1401 -3634 1405 -3630
rect 274 -3810 278 -3806
rect 281 -3810 285 -3806
rect 274 -3817 278 -3813
rect 281 -3817 285 -3813
rect 274 -3824 278 -3820
rect 281 -3824 285 -3820
rect 594 -3810 598 -3806
rect 601 -3810 605 -3806
rect 594 -3817 598 -3813
rect 601 -3817 605 -3813
rect 594 -3824 598 -3820
rect 601 -3824 605 -3820
rect 914 -3810 918 -3806
rect 921 -3810 925 -3806
rect 914 -3817 918 -3813
rect 921 -3817 925 -3813
rect 914 -3824 918 -3820
rect 921 -3824 925 -3820
rect 1234 -3810 1238 -3806
rect 1241 -3810 1245 -3806
rect 1234 -3817 1238 -3813
rect 1241 -3817 1245 -3813
rect 1234 -3824 1238 -3820
rect 1241 -3824 1245 -3820
<< psubstratepdiff >>
rect 118 -3620 121 -3616
rect 114 -3623 125 -3620
rect 118 -3627 121 -3623
rect 114 -3630 125 -3627
rect 118 -3634 121 -3630
rect 438 -3620 441 -3616
rect 434 -3623 445 -3620
rect 438 -3627 441 -3623
rect 434 -3630 445 -3627
rect 438 -3634 441 -3630
rect 758 -3620 761 -3616
rect 754 -3623 765 -3620
rect 758 -3627 761 -3623
rect 754 -3630 765 -3627
rect 758 -3634 761 -3630
rect 1078 -3620 1081 -3616
rect 1074 -3623 1085 -3620
rect 1078 -3627 1081 -3623
rect 1074 -3630 1085 -3627
rect 1078 -3634 1081 -3630
rect 1398 -3620 1401 -3616
rect 1394 -3623 1405 -3620
rect 1398 -3627 1401 -3623
rect 1394 -3630 1405 -3627
rect 1398 -3634 1401 -3630
rect 278 -3810 281 -3806
rect 274 -3813 285 -3810
rect 278 -3817 281 -3813
rect 274 -3820 285 -3817
rect 278 -3824 281 -3820
rect 598 -3810 601 -3806
rect 594 -3813 605 -3810
rect 598 -3817 601 -3813
rect 594 -3820 605 -3817
rect 598 -3824 601 -3820
rect 918 -3810 921 -3806
rect 914 -3813 925 -3810
rect 918 -3817 921 -3813
rect 914 -3820 925 -3817
rect 918 -3824 921 -3820
rect 1238 -3810 1241 -3806
rect 1234 -3813 1245 -3810
rect 1238 -3817 1241 -3813
rect 1234 -3820 1245 -3817
rect 1238 -3824 1241 -3820
<< glass >>
rect 3 -3677 77 -3603
rect 163 -3677 237 -3603
rect 323 -3677 397 -3603
rect 483 -3677 557 -3603
rect 643 -3677 717 -3603
rect 803 -3677 877 -3603
rect 963 -3677 1037 -3603
rect 1123 -3677 1197 -3603
rect 1283 -3677 1357 -3603
rect 1443 -3677 1517 -3603
rect 3 -3837 77 -3763
rect 163 -3837 237 -3763
rect 323 -3837 397 -3763
rect 483 -3837 557 -3763
rect 643 -3837 717 -3763
rect 803 -3837 877 -3763
rect 963 -3837 1037 -3763
rect 1123 -3837 1197 -3763
rect 1283 -3837 1357 -3763
rect 1443 -3837 1517 -3763
<< end >>
