magic
tech scmos
timestamp 617922547
<< ndiffusion >>
rect 0 0 10 3
<< labels >>
rlabel ndiffusion 0 0 0 2 3 B
<< end >>
