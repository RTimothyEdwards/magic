magic
tech scmos
timestamp 616454097
<< polysilicon >>
rect 97 -18 98 -16
rect 106 -18 108 -16
rect 99 -24 101 -22
rect 112 -24 119 -22
rect 122 -24 124 -22
rect 142 -22 149 -20
rect 154 -19 163 -17
rect 142 -24 144 -22
rect 112 -32 114 -24
rect 142 -29 144 -27
rect 106 -36 112 -34
rect 168 -32 170 -30
rect 161 -38 163 -36
rect 171 -38 172 -36
rect 106 -51 114 -50
rect 161 -51 163 -49
rect 171 -51 172 -49
rect 106 -52 112 -51
rect 99 -65 101 -63
rect 112 -63 114 -55
rect 142 -60 144 -58
rect 168 -57 170 -55
rect 112 -65 119 -63
rect 122 -65 124 -63
rect 97 -71 98 -69
rect 106 -71 108 -69
rect 142 -65 144 -63
rect 142 -67 149 -65
rect 154 -70 163 -68
<< ndiffusion >>
rect 98 -14 101 -13
rect 105 -14 106 -13
rect 98 -16 106 -14
rect 163 -14 172 -9
rect 163 -17 173 -14
rect 98 -21 106 -18
rect 102 -24 106 -21
rect 96 -36 99 -24
rect 101 -28 102 -24
rect 101 -34 106 -28
rect 163 -28 168 -19
rect 167 -30 168 -28
rect 170 -30 173 -17
rect 163 -33 167 -32
rect 163 -36 171 -33
rect 96 -39 106 -36
rect 96 -49 97 -39
rect 101 -49 106 -39
rect 163 -41 171 -38
rect 163 -49 171 -46
rect 96 -50 106 -49
rect 96 -63 99 -50
rect 101 -59 106 -52
rect 101 -63 102 -59
rect 102 -66 106 -63
rect 163 -54 171 -51
rect 163 -57 167 -54
rect 167 -61 168 -57
rect 98 -69 106 -66
rect 163 -68 168 -61
rect 170 -70 173 -57
rect 98 -74 106 -71
rect 163 -73 173 -70
rect 163 -75 167 -73
<< pdiffusion >>
rect 119 -21 141 -17
rect 119 -22 122 -21
rect 126 -24 141 -21
rect 119 -25 122 -24
rect 130 -25 137 -24
rect 141 -27 142 -24
rect 144 -27 148 -24
rect 145 -32 148 -27
rect 119 -63 122 -62
rect 130 -63 137 -62
rect 145 -60 148 -55
rect 141 -63 142 -60
rect 144 -63 148 -60
rect 119 -66 122 -65
rect 126 -66 141 -63
rect 119 -70 141 -66
<< metal1 >>
rect 105 -13 107 -9
rect 114 -14 163 -11
rect 90 -19 92 -17
rect 114 -17 117 -14
rect 97 -19 117 -17
rect 90 -20 117 -19
rect 120 -21 149 -17
rect 120 -25 123 -21
rect 160 -21 163 -14
rect 160 -24 177 -21
rect 106 -28 118 -25
rect 122 -29 123 -25
rect 130 -26 137 -24
rect 130 -28 131 -26
rect 136 -28 137 -26
rect 145 -32 163 -29
rect 90 -35 109 -32
rect 106 -39 109 -35
rect 117 -36 144 -33
rect 151 -36 177 -35
rect 151 -38 172 -36
rect 151 -39 154 -38
rect 96 -43 97 -39
rect 92 -44 97 -43
rect 95 -49 97 -44
rect 106 -42 154 -39
rect 106 -48 154 -45
rect 162 -46 165 -41
rect 106 -52 109 -48
rect 151 -49 154 -48
rect 151 -51 172 -49
rect 90 -55 109 -52
rect 117 -54 144 -51
rect 151 -52 177 -51
rect 145 -57 148 -55
rect 106 -62 118 -59
rect 119 -66 122 -62
rect 130 -61 131 -59
rect 136 -61 137 -59
rect 130 -63 137 -61
rect 145 -60 163 -57
rect 90 -68 116 -67
rect 90 -70 92 -68
rect 97 -70 116 -68
rect 119 -70 149 -66
rect 160 -67 177 -64
rect 113 -73 116 -70
rect 160 -73 163 -67
rect 113 -76 163 -73
rect 171 -74 177 -70
rect 171 -78 172 -74
<< metal2 >>
rect 92 -44 97 -9
rect 111 -13 115 -9
rect 110 -14 115 -13
rect 95 -49 97 -44
rect 92 -80 97 -49
rect 111 -80 115 -14
rect 131 -26 136 -9
rect 131 -57 136 -30
rect 131 -80 136 -61
rect 142 -80 146 -9
rect 151 -41 155 -9
rect 151 -46 157 -41
rect 151 -80 155 -46
rect 172 -74 177 -9
rect 172 -80 177 -78
<< polycontact >>
rect 92 -19 97 -14
rect 149 -22 154 -17
rect 112 -36 117 -32
rect 172 -41 177 -36
rect 172 -51 177 -46
rect 112 -55 117 -51
rect 92 -73 97 -68
rect 149 -70 154 -65
<< ndcontact >>
rect 101 -14 105 -9
rect 102 -28 106 -24
rect 163 -32 167 -28
rect 97 -49 101 -39
rect 165 -46 169 -41
rect 102 -63 106 -59
rect 163 -61 167 -57
rect 167 -80 171 -73
<< pdcontact >>
rect 118 -29 122 -25
rect 137 -28 141 -24
rect 144 -36 148 -32
rect 144 -55 148 -51
rect 118 -62 122 -58
rect 137 -63 141 -59
<< m2contact >>
rect 107 -13 111 -9
rect 131 -30 136 -26
rect 91 -49 95 -44
rect 157 -46 162 -41
rect 131 -61 136 -57
rect 172 -78 177 -74
<< ntransistor >>
rect 98 -18 106 -16
rect 99 -34 101 -24
rect 163 -19 170 -17
rect 99 -36 106 -34
rect 168 -30 170 -19
rect 163 -38 171 -36
rect 99 -52 106 -50
rect 163 -51 171 -49
rect 99 -63 101 -52
rect 98 -71 106 -69
rect 168 -68 170 -57
rect 163 -70 170 -68
<< ptransistor >>
rect 119 -24 122 -22
rect 142 -27 144 -24
rect 142 -63 144 -60
rect 119 -65 122 -63
<< psubstratepcontact >>
rect 172 -14 177 -9
rect 92 -43 96 -39
<< nsubstratencontact >>
rect 126 -28 130 -24
rect 126 -63 130 -59
<< labels >>
rlabel metal2 153 -80 153 -80 1 busB0#
rlabel metal2 134 -80 134 -80 1 Vdd!
rlabel metal1 90 -54 90 -54 3 accB1#
rlabel metal1 90 -33 90 -33 3 accB0#
rlabel metal2 113 -80 113 -80 1 busA0#
rlabel metal2 95 -80 95 -80 2 GND!
rlabel metal1 90 -18 90 -18 3 accA0#
rlabel metal1 90 -69 90 -69 3 accA1#
rlabel metal2 174 -80 174 -80 1 GND!
<< end >>
