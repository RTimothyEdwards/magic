magic
tech scmos
timestamp 760840748
<< polysilicon >>
rect 1 87 118 91
rect 1 76 5 87
rect 7 84 13 85
rect 7 80 8 84
rect 12 80 13 84
rect 7 79 13 80
rect 16 84 22 85
rect 16 80 17 84
rect 21 80 22 84
rect 16 79 22 80
rect 25 84 31 85
rect 25 80 26 84
rect 30 80 31 84
rect 25 79 31 80
rect 34 84 40 85
rect 34 80 35 84
rect 39 80 40 84
rect 34 79 40 80
rect 43 84 49 85
rect 43 80 44 84
rect 48 80 49 84
rect 43 79 49 80
rect 52 84 58 85
rect 52 80 53 84
rect 57 80 58 84
rect 52 79 58 80
rect 10 76 13 79
rect 19 76 22 79
rect 28 76 31 79
rect 37 76 40 79
rect 46 76 49 79
rect 1 75 7 76
rect 1 71 2 75
rect 6 71 7 75
rect 10 73 16 76
rect 19 73 25 76
rect 28 73 34 76
rect 37 73 43 76
rect 46 73 52 76
rect 1 70 7 71
rect 13 70 16 73
rect 22 70 25 73
rect 31 70 34 73
rect 40 70 43 73
rect 13 67 19 70
rect 22 67 28 70
rect 31 67 37 70
rect 40 67 46 70
rect 16 64 19 67
rect 25 64 28 67
rect 34 64 37 67
rect 16 61 22 64
rect 25 61 31 64
rect 34 61 40 64
rect 19 58 22 61
rect 28 58 31 61
rect 19 55 25 58
rect 28 55 34 58
rect 22 52 25 55
rect 22 49 28 52
rect 25 -65 28 49
rect 22 -68 28 -65
rect 22 -71 25 -68
rect 31 -71 34 55
rect 19 -74 25 -71
rect 28 -74 34 -71
rect 19 -77 22 -74
rect 28 -77 31 -74
rect 37 -77 40 61
rect 16 -80 22 -77
rect 25 -80 31 -77
rect 34 -80 40 -77
rect 16 -95 19 -80
rect 25 -95 28 -80
rect 34 -95 37 -80
rect 43 -95 46 67
rect 49 -89 52 73
rect 55 -83 58 79
rect 61 84 67 85
rect 61 80 62 84
rect 66 80 67 84
rect 61 79 67 80
rect 70 84 76 85
rect 70 80 71 84
rect 75 80 76 84
rect 70 79 76 80
rect 79 84 85 85
rect 79 80 80 84
rect 84 80 85 84
rect 79 79 85 80
rect 88 84 94 85
rect 88 80 89 84
rect 93 80 94 84
rect 88 79 94 80
rect 97 84 103 85
rect 97 80 98 84
rect 102 80 103 84
rect 97 79 103 80
rect 106 84 112 85
rect 106 80 107 84
rect 111 80 112 84
rect 106 79 112 80
rect 61 -77 64 79
rect 70 76 73 79
rect 79 76 82 79
rect 88 76 91 79
rect 97 76 100 79
rect 106 76 109 79
rect 114 76 118 87
rect 67 73 73 76
rect 76 73 82 76
rect 85 73 91 76
rect 94 73 100 76
rect 103 73 109 76
rect 112 75 118 76
rect 67 -71 70 73
rect 76 70 79 73
rect 85 70 88 73
rect 94 70 97 73
rect 103 70 106 73
rect 112 71 113 75
rect 117 71 118 75
rect 112 70 118 71
rect 73 67 79 70
rect 82 67 88 70
rect 91 67 97 70
rect 100 67 106 70
rect 73 -65 76 67
rect 82 64 85 67
rect 91 64 94 67
rect 100 64 103 67
rect 79 61 85 64
rect 88 61 94 64
rect 97 61 103 64
rect 79 -59 82 61
rect 88 58 91 61
rect 97 58 100 61
rect 85 55 91 58
rect 94 55 100 58
rect 85 -53 88 55
rect 94 52 97 55
rect 91 49 97 52
rect 91 -47 94 49
rect 91 -50 100 -47
rect 85 -56 94 -53
rect 79 -62 88 -59
rect 73 -68 82 -65
rect 67 -74 76 -71
rect 61 -80 70 -77
rect 55 -86 64 -83
rect 49 -92 55 -89
rect 52 -95 55 -92
rect 61 -95 64 -86
rect 67 -89 70 -80
rect 73 -83 76 -74
rect 79 -77 82 -68
rect 85 -71 88 -62
rect 91 -65 94 -56
rect 97 -59 100 -50
rect 97 -62 103 -59
rect 100 -65 103 -62
rect 91 -68 97 -65
rect 100 -68 106 -65
rect 94 -71 97 -68
rect 103 -71 106 -68
rect 85 -74 91 -71
rect 94 -74 100 -71
rect 103 -74 109 -71
rect 88 -77 91 -74
rect 97 -77 100 -74
rect 106 -77 109 -74
rect 79 -80 85 -77
rect 88 -80 94 -77
rect 97 -80 103 -77
rect 106 -80 112 -77
rect 82 -83 85 -80
rect 91 -83 94 -80
rect 100 -83 103 -80
rect 109 -83 112 -80
rect 73 -86 79 -83
rect 82 -86 88 -83
rect 91 -86 97 -83
rect 100 -86 106 -83
rect 109 -86 115 -83
rect 76 -89 79 -86
rect 85 -89 88 -86
rect 94 -89 97 -86
rect 103 -89 106 -86
rect 112 -88 115 -86
rect 67 -92 73 -89
rect 76 -92 82 -89
rect 85 -92 91 -89
rect 94 -92 100 -89
rect 103 -92 109 -89
rect 112 -91 118 -88
rect 70 -95 73 -92
rect 79 -95 82 -92
rect 88 -95 91 -92
rect 97 -95 100 -92
rect 106 -95 109 -92
rect 115 -95 118 -91
rect 16 -96 22 -95
rect 16 -100 17 -96
rect 21 -100 22 -96
rect 16 -101 22 -100
rect 25 -96 31 -95
rect 25 -100 26 -96
rect 30 -100 31 -96
rect 25 -101 31 -100
rect 34 -96 40 -95
rect 34 -100 35 -96
rect 39 -100 40 -96
rect 34 -101 40 -100
rect 43 -96 49 -95
rect 43 -100 44 -96
rect 48 -100 49 -96
rect 43 -101 49 -100
rect 52 -96 58 -95
rect 52 -100 53 -96
rect 57 -100 58 -96
rect 52 -101 58 -100
rect 61 -96 67 -95
rect 61 -100 62 -96
rect 66 -100 67 -96
rect 61 -101 67 -100
rect 70 -96 76 -95
rect 70 -100 71 -96
rect 75 -100 76 -96
rect 70 -101 76 -100
rect 79 -96 85 -95
rect 79 -100 80 -96
rect 84 -100 85 -96
rect 79 -101 85 -100
rect 88 -96 94 -95
rect 88 -100 89 -96
rect 93 -100 94 -96
rect 88 -101 94 -100
rect 97 -96 103 -95
rect 97 -100 98 -96
rect 102 -100 103 -96
rect 97 -101 103 -100
rect 106 -96 112 -95
rect 106 -100 107 -96
rect 111 -100 112 -96
rect 106 -101 112 -100
rect 115 -96 121 -95
rect 115 -100 116 -96
rect 120 -100 121 -96
rect 115 -101 121 -100
<< metal1 >>
rect 7 84 13 85
rect 7 80 8 84
rect 12 80 13 84
rect 7 79 13 80
rect 16 84 22 85
rect 16 80 17 84
rect 21 80 22 84
rect 16 79 22 80
rect 25 84 31 85
rect 25 80 26 84
rect 30 80 31 84
rect 25 79 31 80
rect 34 84 40 85
rect 34 80 35 84
rect 39 80 40 84
rect 34 79 40 80
rect 43 84 49 85
rect 43 80 44 84
rect 48 80 49 84
rect 43 79 49 80
rect 52 84 58 85
rect 52 80 53 84
rect 57 80 58 84
rect 52 79 58 80
rect 10 76 13 79
rect 19 76 22 79
rect 28 76 31 79
rect 37 76 40 79
rect 46 76 49 79
rect 1 75 7 76
rect 1 71 2 75
rect 6 71 7 75
rect 10 73 16 76
rect 19 73 25 76
rect 28 73 34 76
rect 37 73 43 76
rect 46 73 52 76
rect 1 70 7 71
rect 13 70 16 73
rect 22 70 25 73
rect 31 70 34 73
rect 40 70 43 73
rect 4 67 10 70
rect 13 67 19 70
rect 22 67 28 70
rect 31 67 37 70
rect 40 67 46 70
rect 7 64 10 67
rect 16 64 19 67
rect 25 64 28 67
rect 34 64 37 67
rect 7 61 13 64
rect 16 61 22 64
rect 25 61 31 64
rect 34 61 40 64
rect 10 58 13 61
rect 19 58 22 61
rect 28 58 31 61
rect 10 55 16 58
rect 19 55 25 58
rect 28 55 34 58
rect 13 52 16 55
rect 22 52 25 55
rect 13 49 19 52
rect 22 49 28 52
rect 16 46 19 49
rect 16 43 22 46
rect 19 -59 22 43
rect 16 -62 22 -59
rect 16 -65 19 -62
rect 25 -65 28 49
rect 13 -68 19 -65
rect 22 -68 28 -65
rect 13 -71 16 -68
rect 22 -71 25 -68
rect 31 -71 34 55
rect 10 -74 16 -71
rect 19 -74 25 -71
rect 28 -74 34 -71
rect 10 -77 13 -74
rect 19 -77 22 -74
rect 28 -77 31 -74
rect 37 -77 40 61
rect 4 -80 13 -77
rect 16 -80 22 -77
rect 25 -80 31 -77
rect 34 -80 40 -77
rect 4 -110 7 -80
rect 16 -83 19 -80
rect 25 -83 28 -80
rect 34 -83 37 -80
rect 43 -83 46 67
rect 10 -86 19 -83
rect 22 -86 28 -83
rect 31 -86 37 -83
rect 40 -86 46 -83
rect 10 -110 13 -86
rect 22 -89 25 -86
rect 31 -89 34 -86
rect 40 -89 43 -86
rect 49 -89 52 73
rect 19 -92 25 -89
rect 28 -92 34 -89
rect 37 -92 43 -89
rect 46 -92 52 -89
rect 19 -95 22 -92
rect 28 -95 31 -92
rect 37 -95 40 -92
rect 46 -95 49 -92
rect 55 -95 58 79
rect 16 -96 22 -95
rect 16 -100 17 -96
rect 21 -100 22 -96
rect 16 -101 22 -100
rect 25 -96 31 -95
rect 25 -100 26 -96
rect 30 -100 31 -96
rect 25 -101 31 -100
rect 34 -96 40 -95
rect 34 -100 35 -96
rect 39 -100 40 -96
rect 34 -101 40 -100
rect 43 -96 49 -95
rect 43 -100 44 -96
rect 48 -100 49 -96
rect 43 -101 49 -100
rect 52 -96 58 -95
rect 52 -100 53 -96
rect 57 -100 58 -96
rect 52 -101 58 -100
rect 61 84 67 85
rect 61 80 62 84
rect 66 80 67 84
rect 61 79 67 80
rect 70 84 76 85
rect 70 80 71 84
rect 75 80 76 84
rect 70 79 76 80
rect 79 84 85 85
rect 79 80 80 84
rect 84 80 85 84
rect 79 79 85 80
rect 88 84 94 85
rect 88 80 89 84
rect 93 80 94 84
rect 88 79 94 80
rect 97 84 103 85
rect 97 80 98 84
rect 102 80 103 84
rect 97 79 103 80
rect 106 84 112 85
rect 106 80 107 84
rect 111 80 112 84
rect 106 79 112 80
rect 61 -95 64 79
rect 70 76 73 79
rect 79 76 82 79
rect 88 76 91 79
rect 97 76 100 79
rect 106 76 109 79
rect 67 73 73 76
rect 76 73 82 76
rect 85 73 91 76
rect 94 73 100 76
rect 103 73 109 76
rect 112 75 118 76
rect 67 -89 70 73
rect 76 70 79 73
rect 85 70 88 73
rect 94 70 97 73
rect 103 70 106 73
rect 112 71 113 75
rect 117 71 118 75
rect 112 70 118 71
rect 73 67 79 70
rect 82 67 88 70
rect 91 67 97 70
rect 100 67 106 70
rect 109 67 115 70
rect 73 -83 76 67
rect 82 64 85 67
rect 91 64 94 67
rect 100 64 103 67
rect 109 64 112 67
rect 79 61 85 64
rect 88 61 94 64
rect 97 61 103 64
rect 106 61 112 64
rect 79 -77 82 61
rect 88 58 91 61
rect 97 58 100 61
rect 106 58 109 61
rect 85 55 91 58
rect 94 55 100 58
rect 103 55 109 58
rect 85 -71 88 55
rect 94 52 97 55
rect 103 52 106 55
rect 91 49 97 52
rect 100 49 106 52
rect 91 -65 94 49
rect 100 46 103 49
rect 97 43 103 46
rect 97 -59 100 43
rect 97 -62 103 -59
rect 100 -65 103 -62
rect 91 -68 97 -65
rect 100 -68 106 -65
rect 94 -71 97 -68
rect 103 -71 106 -68
rect 85 -74 91 -71
rect 94 -74 100 -71
rect 103 -74 109 -71
rect 88 -77 91 -74
rect 97 -77 100 -74
rect 106 -77 109 -74
rect 79 -80 85 -77
rect 88 -80 94 -77
rect 97 -80 103 -77
rect 106 -80 112 -77
rect 82 -83 85 -80
rect 91 -83 94 -80
rect 100 -83 103 -80
rect 109 -83 112 -80
rect 73 -86 79 -83
rect 82 -86 88 -83
rect 91 -86 97 -83
rect 100 -86 106 -83
rect 109 -86 115 -83
rect 76 -89 79 -86
rect 85 -89 88 -86
rect 94 -89 97 -86
rect 103 -89 106 -86
rect 112 -88 115 -86
rect 67 -92 73 -89
rect 76 -92 82 -89
rect 85 -92 91 -89
rect 94 -92 100 -89
rect 103 -92 109 -89
rect 112 -91 127 -88
rect 70 -95 73 -92
rect 79 -95 82 -92
rect 88 -95 91 -92
rect 97 -95 100 -92
rect 106 -95 109 -92
rect 61 -96 67 -95
rect 61 -100 62 -96
rect 66 -100 67 -96
rect 61 -101 67 -100
rect 70 -96 76 -95
rect 70 -100 71 -96
rect 75 -100 76 -96
rect 70 -101 76 -100
rect 79 -96 85 -95
rect 79 -100 80 -96
rect 84 -100 85 -96
rect 79 -101 85 -100
rect 88 -96 94 -95
rect 88 -100 89 -96
rect 93 -100 94 -96
rect 88 -101 94 -100
rect 97 -96 103 -95
rect 97 -100 98 -96
rect 102 -100 103 -96
rect 97 -101 103 -100
rect 106 -96 112 -95
rect 106 -100 107 -96
rect 111 -100 112 -96
rect 106 -101 112 -100
rect 115 -96 121 -95
rect 115 -100 116 -96
rect 120 -100 121 -96
rect 115 -101 121 -100
rect 115 -110 118 -101
rect 124 -110 127 -91
<< polycontact >>
rect 8 80 12 84
rect 17 80 21 84
rect 26 80 30 84
rect 35 80 39 84
rect 44 80 48 84
rect 53 80 57 84
rect 2 71 6 75
rect 62 80 66 84
rect 71 80 75 84
rect 80 80 84 84
rect 89 80 93 84
rect 98 80 102 84
rect 107 80 111 84
rect 113 71 117 75
rect 17 -100 21 -96
rect 26 -100 30 -96
rect 35 -100 39 -96
rect 44 -100 48 -96
rect 53 -100 57 -96
rect 62 -100 66 -96
rect 71 -100 75 -96
rect 80 -100 84 -96
rect 89 -100 93 -96
rect 98 -100 102 -96
rect 107 -100 111 -96
rect 116 -100 120 -96
<< substrateopen >>
rect -16 94 134 110
rect -16 67 -3 94
rect 121 67 134 94
rect -16 64 0 67
rect 118 64 134 67
rect -16 58 3 64
rect 115 58 134 64
rect -16 52 6 58
rect 112 52 134 58
rect -16 46 9 52
rect 109 46 134 52
rect -16 40 12 46
rect 106 40 134 46
rect -16 -10 16 40
rect 102 -10 134 40
<< labels >>
rlabel metal1 125 -109 125 -109 8 heater2
rlabel metal1 5 -109 5 -109 8 heater1
rlabel metal1 11 -109 11 -109 8 Vmeas1
rlabel metal1 116 -109 116 -109 8 Vmeas2
<< end >>
