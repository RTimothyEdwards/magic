magic
tech scmos
timestamp 760840453
<< substrateopen >>
rect 647 -163 707 -162
rect 648 -164 706 -163
rect 649 -165 705 -164
rect 650 -166 704 -165
rect 651 -167 703 -166
rect 652 -168 702 -167
rect 653 -169 701 -168
rect 654 -170 700 -169
rect 655 -171 699 -170
rect 656 -172 698 -171
rect 637 -173 638 -172
rect 657 -173 697 -172
rect 716 -173 717 -172
rect 637 -174 639 -173
rect 658 -174 696 -173
rect 715 -174 717 -173
rect 637 -175 640 -174
rect 659 -175 695 -174
rect 714 -175 717 -174
rect 637 -176 641 -175
rect 660 -176 694 -175
rect 713 -176 717 -175
rect 637 -177 642 -176
rect 661 -177 693 -176
rect 712 -177 717 -176
rect 637 -178 643 -177
rect 662 -178 692 -177
rect 711 -178 717 -177
rect 637 -179 644 -178
rect 663 -179 691 -178
rect 710 -179 717 -178
rect 637 -180 645 -179
rect 664 -180 690 -179
rect 709 -180 717 -179
rect 637 -181 646 -180
rect 665 -181 689 -180
rect 708 -181 717 -180
rect 637 -182 647 -181
rect 707 -182 717 -181
rect 637 -183 648 -182
rect 706 -183 717 -182
rect 637 -184 649 -183
rect 705 -184 717 -183
rect 637 -185 650 -184
rect 704 -185 717 -184
rect 637 -186 651 -185
rect 703 -186 717 -185
rect 637 -187 652 -186
rect 702 -187 717 -186
rect 637 -188 653 -187
rect 701 -188 717 -187
rect 637 -189 654 -188
rect 700 -189 717 -188
rect 637 -190 655 -189
rect 699 -190 717 -189
rect 637 -214 656 -190
rect 698 -214 717 -190
rect 637 -215 655 -214
rect 699 -215 717 -214
rect 637 -216 654 -215
rect 700 -216 717 -215
rect 637 -217 653 -216
rect 701 -217 717 -216
rect 637 -218 652 -217
rect 702 -218 717 -217
rect 637 -219 651 -218
rect 703 -219 717 -218
rect 637 -220 650 -219
rect 704 -220 717 -219
rect 637 -221 649 -220
rect 705 -221 717 -220
rect 637 -222 648 -221
rect 706 -222 717 -221
rect 637 -223 647 -222
rect 707 -223 717 -222
rect 637 -224 646 -223
rect 665 -224 689 -223
rect 708 -224 717 -223
rect 637 -225 645 -224
rect 664 -225 690 -224
rect 709 -225 717 -224
rect 637 -226 644 -225
rect 663 -226 691 -225
rect 710 -226 717 -225
rect 637 -227 643 -226
rect 662 -227 692 -226
rect 711 -227 717 -226
rect 637 -228 642 -227
rect 661 -228 693 -227
rect 712 -228 717 -227
rect 637 -229 641 -228
rect 660 -229 694 -228
rect 713 -229 717 -228
rect 637 -230 640 -229
rect 659 -230 695 -229
rect 714 -230 717 -229
rect 637 -231 639 -230
rect 658 -231 696 -230
rect 715 -231 717 -230
rect 637 -232 638 -231
rect 657 -232 697 -231
rect 716 -232 717 -231
rect 656 -233 698 -232
rect 655 -234 699 -233
rect 654 -235 700 -234
rect 653 -236 701 -235
rect 652 -237 702 -236
rect 651 -238 703 -237
rect 650 -239 704 -238
rect 649 -240 705 -239
rect 648 -241 706 -240
rect 647 -242 707 -241
<< end >>
