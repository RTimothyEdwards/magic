magic
tech scmos
timestamp 801255023
<< nwell >>
rect -4 52 96 140
rect 0 -2 92 43
<< metal1 >>
rect 21 124 39 128
rect 65 124 83 128
rect 10 110 28 114
rect 54 110 72 114
rect -5 75 17 79
rect 43 75 61 79
rect 83 65 87 75
rect -5 61 6 65
rect 32 61 50 65
rect 76 61 87 65
rect 78 34 92 35
rect 78 30 79 34
rect 83 30 92 34
rect 78 29 92 30
rect 0 11 14 12
rect 0 7 9 11
rect 13 7 14 11
rect 0 6 14 7
<< pbase >>
rect 14 128 24 131
rect 14 124 17 128
rect 21 124 24 128
rect 14 121 24 124
rect 36 128 46 131
rect 36 124 39 128
rect 43 124 46 128
rect 36 121 46 124
rect 58 128 68 131
rect 58 124 61 128
rect 65 124 68 128
rect 58 121 68 124
rect 80 128 90 131
rect 80 124 83 128
rect 87 124 90 128
rect 80 121 90 124
rect 3 114 13 117
rect 3 110 6 114
rect 10 110 13 114
rect 3 107 13 110
rect 6 68 10 107
rect 17 82 21 121
rect 25 114 35 117
rect 25 110 28 114
rect 32 110 35 114
rect 25 107 35 110
rect 14 79 24 82
rect 14 75 17 79
rect 21 75 24 79
rect 14 72 24 75
rect 28 68 32 107
rect 39 82 43 121
rect 47 114 57 117
rect 47 110 50 114
rect 54 110 57 114
rect 47 107 57 110
rect 36 79 46 82
rect 36 75 39 79
rect 43 75 46 79
rect 36 72 46 75
rect 50 68 54 107
rect 61 82 65 121
rect 69 114 79 117
rect 69 110 72 114
rect 76 110 79 114
rect 69 107 79 110
rect 58 79 68 82
rect 58 75 61 79
rect 65 75 68 79
rect 58 72 68 75
rect 72 68 76 107
rect 83 82 87 121
rect 80 79 90 82
rect 80 75 83 79
rect 87 75 90 79
rect 80 72 90 75
rect 3 65 13 68
rect 3 61 6 65
rect 10 61 13 65
rect 3 58 13 61
rect 25 65 35 68
rect 25 61 28 65
rect 32 61 35 65
rect 25 58 35 61
rect 47 65 57 68
rect 47 61 50 65
rect 54 61 57 65
rect 47 58 57 61
rect 69 65 79 68
rect 69 61 72 65
rect 76 61 79 65
rect 69 58 79 61
rect 9 33 24 37
rect 9 14 13 33
rect 6 11 16 14
rect 6 7 9 11
rect 13 7 16 11
rect 6 4 16 7
rect 20 8 24 33
rect 28 33 40 37
rect 28 8 32 33
rect 20 4 32 8
rect 36 8 40 33
rect 44 33 56 37
rect 44 8 48 33
rect 36 4 48 8
rect 52 8 56 33
rect 60 33 72 37
rect 60 8 64 33
rect 52 4 64 8
rect 68 8 72 33
rect 76 34 86 37
rect 76 30 79 34
rect 83 30 86 34
rect 76 27 86 30
rect 79 8 83 27
rect 68 4 83 8
<< pbasecontact >>
rect 17 124 21 128
rect 39 124 43 128
rect 61 124 65 128
rect 83 124 87 128
rect 6 110 10 114
rect 28 110 32 114
rect 17 75 21 79
rect 50 110 54 114
rect 39 75 43 79
rect 72 110 76 114
rect 61 75 65 79
rect 83 75 87 79
rect 6 61 10 65
rect 28 61 32 65
rect 50 61 54 65
rect 72 61 76 65
rect 9 7 13 11
rect 79 30 83 34
<< labels >>
rlabel metal1 2 9 2 9 3 a
rlabel metal1 90 32 90 32 7 b
<< end >>
