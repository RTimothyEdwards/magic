magic
tech scmos
timestamp 500619087
<< polysilicon >>
rect -6 5 0 7
rect 3 5 10 7
<< ndiffusion >>
rect 0 7 3 8
rect 0 4 3 5
<< metal1 >>
rect -6 8 0 12
rect 4 8 10 12
rect -6 0 0 4
rect 4 0 10 4
<< ndcontact >>
rect 0 8 4 12
rect 0 0 4 4
<< ntransistor >>
rect 0 5 3 7
use tut8d tut8d_0
timestamp 500619087
transform 1 0 0 0 1 3
box 10 -3 18 9
<< labels >>
rlabel metal1 -6 0 -6 4 3 Out
rlabel metal1 -6 8 -6 12 3 In
rlabel polysilicon -6 5 -6 7 3 Gate
<< end >>
