magic
tech scmos
timestamp 783737922
<< nwell >>
rect 18 19 174 135
<< metal1 >>
rect 0 146 179 155
rect 15 139 17 143
rect 44 125 53 127
rect 57 118 63 146
rect 67 125 76 127
rect 116 125 125 127
rect 129 118 135 146
rect 175 139 177 143
rect 139 125 148 127
rect 21 114 35 118
rect 50 114 70 118
rect 85 114 107 118
rect 122 114 142 118
rect 157 114 171 118
rect 21 92 27 114
rect 44 105 53 107
rect 57 92 63 114
rect 67 105 76 107
rect 93 92 99 114
rect 116 105 125 107
rect 129 92 135 114
rect 139 105 148 107
rect 165 92 171 114
rect 21 88 35 92
rect 50 88 70 92
rect 85 88 107 92
rect 122 88 142 92
rect 157 88 171 92
rect 21 66 27 88
rect 44 79 53 81
rect 57 66 63 88
rect 67 79 76 81
rect 93 66 99 88
rect 116 79 125 81
rect 129 66 135 88
rect 139 79 148 81
rect 165 66 171 88
rect 21 62 35 66
rect 50 62 70 66
rect 85 62 107 66
rect 122 62 142 66
rect 157 62 171 66
rect 21 40 27 62
rect 44 53 53 55
rect 57 40 63 62
rect 67 53 76 55
rect 93 40 99 62
rect 116 53 125 55
rect 129 40 135 62
rect 139 53 148 55
rect 165 40 171 62
rect 21 36 35 40
rect 50 36 70 40
rect 85 36 107 40
rect 122 36 142 40
rect 157 36 171 40
rect 21 8 27 36
rect 44 27 53 29
rect 67 27 76 29
rect 93 8 99 36
rect 116 27 125 29
rect 139 27 148 29
rect 165 8 171 36
rect 181 16 182 143
rect 177 15 182 16
rect 180 11 182 15
rect 0 -1 180 8
<< metal2 >>
rect 53 139 68 143
rect 124 139 139 143
rect 175 139 182 143
rect -2 125 149 126
rect -2 121 44 125
rect 53 121 67 125
rect 76 121 116 125
rect 125 121 139 125
rect 148 121 149 125
rect -2 120 149 121
rect -2 112 8 120
rect -2 111 149 112
rect -2 107 44 111
rect 53 107 67 111
rect 76 107 116 111
rect 125 107 139 111
rect 148 107 149 111
rect -2 106 149 107
rect -2 86 8 106
rect -2 85 149 86
rect -2 81 44 85
rect 53 81 67 85
rect 76 81 116 85
rect 125 81 139 85
rect 148 81 149 85
rect -2 80 149 81
rect -2 60 8 80
rect -2 59 59 60
rect -2 55 44 59
rect 53 55 59 59
rect -2 54 59 55
rect 63 59 149 60
rect 63 55 67 59
rect 76 55 116 59
rect 125 55 139 59
rect 148 55 149 59
rect 63 54 149 55
rect -2 34 8 54
rect -2 33 149 34
rect -2 29 44 33
rect 53 29 67 33
rect 76 29 116 33
rect 125 29 139 33
rect 148 29 149 33
rect -2 28 149 29
rect -2 12 8 28
rect 177 15 182 139
rect 90 11 102 15
rect 162 11 176 15
rect 180 11 182 15
rect 186 11 187 143
<< collector >>
rect 21 131 171 132
rect 21 127 22 131
rect 54 127 66 131
rect 126 127 138 131
rect 170 127 171 131
rect 21 126 171 127
rect 21 106 27 126
rect 57 106 63 126
rect 93 106 99 126
rect 129 106 135 126
rect 165 106 171 126
rect 21 105 171 106
rect 21 101 30 105
rect 54 101 66 105
rect 90 101 102 105
rect 126 101 138 105
rect 162 101 171 105
rect 21 100 171 101
rect 21 80 27 100
rect 57 80 63 100
rect 93 80 99 100
rect 129 80 135 100
rect 165 80 171 100
rect 21 79 171 80
rect 21 75 30 79
rect 54 75 66 79
rect 90 75 102 79
rect 126 75 138 79
rect 162 75 171 79
rect 21 74 171 75
rect 21 54 27 74
rect 57 54 63 74
rect 93 54 99 74
rect 129 54 135 74
rect 165 54 171 74
rect 21 53 171 54
rect 21 49 30 53
rect 54 49 66 53
rect 90 49 102 53
rect 126 49 138 53
rect 162 49 171 53
rect 21 48 171 49
rect 21 28 27 48
rect 57 28 63 48
rect 93 28 99 48
rect 129 28 135 48
rect 165 28 171 48
rect 21 27 171 28
rect 21 23 30 27
rect 90 23 102 27
rect 162 23 171 27
rect 21 22 171 23
<< pbase >>
rect 31 118 53 122
rect 31 114 35 118
rect 39 114 46 118
rect 50 114 53 118
rect 31 110 53 114
rect 67 118 89 122
rect 67 114 70 118
rect 74 114 81 118
rect 85 114 89 118
rect 67 110 89 114
rect 103 118 125 122
rect 103 114 107 118
rect 111 114 118 118
rect 122 114 125 118
rect 103 110 125 114
rect 139 118 161 122
rect 139 114 142 118
rect 146 114 153 118
rect 157 114 161 118
rect 139 110 161 114
rect 31 92 53 96
rect 31 88 35 92
rect 39 88 46 92
rect 50 88 53 92
rect 31 84 53 88
rect 67 92 89 96
rect 67 88 70 92
rect 74 88 81 92
rect 85 88 89 92
rect 67 84 89 88
rect 103 92 125 96
rect 103 88 107 92
rect 111 88 118 92
rect 122 88 125 92
rect 103 84 125 88
rect 139 92 161 96
rect 139 88 142 92
rect 146 88 153 92
rect 157 88 161 92
rect 139 84 161 88
rect 31 66 53 70
rect 31 62 35 66
rect 39 62 46 66
rect 50 62 53 66
rect 31 58 53 62
rect 67 66 89 70
rect 67 62 70 66
rect 74 62 81 66
rect 85 62 89 66
rect 67 58 89 62
rect 103 66 125 70
rect 103 62 107 66
rect 111 62 118 66
rect 122 62 125 66
rect 103 58 125 62
rect 139 66 161 70
rect 139 62 142 66
rect 146 62 153 66
rect 157 62 161 66
rect 139 58 161 62
rect 31 40 53 44
rect 31 36 35 40
rect 39 36 46 40
rect 50 36 53 40
rect 31 32 53 36
rect 67 40 89 44
rect 67 36 70 40
rect 74 36 81 40
rect 85 36 89 40
rect 67 32 89 36
rect 103 40 125 44
rect 103 36 107 40
rect 111 36 118 40
rect 122 36 125 40
rect 103 32 125 36
rect 139 40 161 44
rect 139 36 142 40
rect 146 36 153 40
rect 157 36 161 40
rect 139 32 161 36
<< collectorcontact >>
rect 22 127 54 131
rect 66 127 126 131
rect 138 127 170 131
rect 30 101 54 105
rect 66 101 90 105
rect 102 101 126 105
rect 138 101 162 105
rect 30 75 54 79
rect 66 75 90 79
rect 102 75 126 79
rect 138 75 162 79
rect 30 49 54 53
rect 66 49 90 53
rect 102 49 126 53
rect 138 49 162 53
rect 30 23 90 27
rect 102 23 162 27
<< emittercontact >>
rect 35 114 39 118
rect 81 114 85 118
rect 107 114 111 118
rect 153 114 157 118
rect 35 88 39 92
rect 81 88 85 92
rect 107 88 111 92
rect 153 88 157 92
rect 35 62 39 66
rect 81 62 85 66
rect 107 62 111 66
rect 153 62 157 66
rect 35 36 39 40
rect 81 36 85 40
rect 107 36 111 40
rect 153 36 157 40
<< pbasecontact >>
rect 46 114 50 118
rect 70 114 74 118
rect 118 114 122 118
rect 142 114 146 118
rect 46 88 50 92
rect 70 88 74 92
rect 118 88 122 92
rect 142 88 146 92
rect 46 62 50 66
rect 70 62 74 66
rect 118 62 122 66
rect 142 62 146 66
rect 46 36 50 40
rect 70 36 74 40
rect 118 36 122 40
rect 142 36 146 40
<< m2contact >>
rect 17 139 21 143
rect 25 139 29 143
rect 33 139 37 143
rect 41 139 45 143
rect 49 139 53 143
rect 44 121 53 125
rect 68 139 72 143
rect 76 139 80 143
rect 84 139 88 143
rect 92 139 96 143
rect 100 139 104 143
rect 108 139 112 143
rect 116 139 120 143
rect 67 121 76 125
rect 116 121 125 125
rect 139 139 143 143
rect 147 139 151 143
rect 155 139 159 143
rect 163 139 167 143
rect 171 139 175 143
rect 139 121 148 125
rect 44 107 53 111
rect 67 107 76 111
rect 116 107 125 111
rect 139 107 148 111
rect 44 81 53 85
rect 67 81 76 85
rect 116 81 125 85
rect 139 81 148 85
rect 44 55 53 59
rect 67 55 76 59
rect 116 55 125 59
rect 139 55 148 59
rect 44 29 53 33
rect 67 29 76 33
rect 30 11 34 15
rect 38 11 42 15
rect 46 11 50 15
rect 54 11 58 15
rect 62 11 66 15
rect 70 11 74 15
rect 78 11 82 15
rect 86 11 90 15
rect 116 29 125 33
rect 139 29 148 33
rect 102 11 106 15
rect 110 11 114 15
rect 118 11 122 15
rect 126 11 130 15
rect 134 11 138 15
rect 142 11 146 15
rect 150 11 154 15
rect 158 11 162 15
rect 176 11 180 15
rect 182 11 186 143
<< psubstratepcontact >>
rect 11 12 15 143
rect 21 139 25 143
rect 29 139 33 143
rect 37 139 41 143
rect 45 139 49 143
rect 72 139 76 143
rect 80 139 84 143
rect 88 139 92 143
rect 96 139 100 143
rect 104 139 108 143
rect 112 139 116 143
rect 120 139 124 143
rect 143 139 147 143
rect 151 139 155 143
rect 159 139 163 143
rect 167 139 171 143
rect 177 16 181 143
rect 34 11 38 15
rect 42 11 46 15
rect 50 11 54 15
rect 58 11 62 15
rect 66 11 70 15
rect 74 11 78 15
rect 82 11 86 15
rect 106 11 110 15
rect 114 11 118 15
rect 122 11 126 15
rect 130 11 134 15
rect 138 11 142 15
rect 146 11 150 15
rect 154 11 158 15
<< psubstratepdiff >>
rect 11 143 181 144
rect 15 139 21 143
rect 25 139 29 143
rect 33 139 37 143
rect 41 139 45 143
rect 49 139 72 143
rect 76 139 80 143
rect 84 139 88 143
rect 92 139 96 143
rect 100 139 104 143
rect 108 139 112 143
rect 116 139 120 143
rect 124 139 143 143
rect 147 139 151 143
rect 155 139 159 143
rect 163 139 167 143
rect 171 139 177 143
rect 15 138 177 139
rect 15 15 181 16
rect 15 12 34 15
rect 11 11 34 12
rect 38 11 42 15
rect 46 11 50 15
rect 54 11 58 15
rect 62 11 66 15
rect 70 11 74 15
rect 78 11 82 15
rect 86 11 106 15
rect 110 11 114 15
rect 118 11 122 15
rect 126 11 130 15
rect 134 11 138 15
rect 142 11 146 15
rect 150 11 154 15
rect 158 11 181 15
rect 11 10 181 11
<< labels >>
rlabel metal1 0 -1 179 8 0 emitter
rlabel metal2 187 13 187 140 7 GND
rlabel metal1 0 146 179 155 0 base
rlabel metal2 -2 13 8 125 0 collector
<< end >>
