magic
tech scmos
timestamp 765071885
<< polysilicon >>
rect 72 492 92 493
rect 71 491 92 492
rect 70 490 93 491
rect 69 489 93 490
rect 68 488 94 489
rect 67 487 94 488
rect 66 486 95 487
rect 65 485 95 486
rect 64 484 96 485
rect 63 483 96 484
rect 62 482 97 483
rect 61 481 97 482
rect 60 480 98 481
rect 59 479 98 480
rect 58 478 99 479
rect 57 477 99 478
rect 56 476 100 477
rect 55 475 100 476
rect 54 474 101 475
rect 53 473 101 474
rect 52 471 102 473
rect 52 469 103 471
rect 52 467 104 469
rect 52 465 105 467
rect 52 463 106 465
rect 52 461 107 463
rect 52 460 108 461
rect 52 459 78 460
rect 79 459 108 460
rect 52 458 77 459
rect 52 457 76 458
rect 80 457 109 459
rect 52 456 75 457
rect 52 455 74 456
rect 81 455 110 457
rect 52 454 73 455
rect 52 313 72 454
rect 82 453 111 455
rect 83 451 112 453
rect 84 449 113 451
rect 85 447 114 449
rect 86 445 115 447
rect 87 443 116 445
rect 88 441 117 443
rect 89 439 118 441
rect 90 437 119 439
rect 91 435 120 437
rect 92 433 121 435
rect 93 431 122 433
rect 94 429 123 431
rect 95 427 124 429
rect 96 425 125 427
rect 97 423 126 425
rect 98 421 127 423
rect 99 419 128 421
rect 100 417 129 419
rect 101 415 130 417
rect 102 413 131 415
rect 103 411 132 413
rect 104 409 133 411
rect 105 407 134 409
rect 106 405 135 407
rect 107 403 136 405
rect 108 401 137 403
rect 109 399 138 401
rect 110 397 139 399
rect 111 395 140 397
rect 112 393 141 395
rect 113 391 142 393
rect 114 389 143 391
rect 115 387 144 389
rect 116 385 145 387
rect 117 383 146 385
rect 118 381 147 383
rect 119 379 148 381
rect 120 377 149 379
rect 121 375 150 377
rect 122 373 151 375
rect 123 371 152 373
rect 124 369 153 371
rect 125 367 154 369
rect 126 365 155 367
rect 127 363 156 365
rect 128 361 157 363
rect 129 359 158 361
rect 130 357 159 359
rect 131 355 160 357
rect 132 353 161 355
rect 133 351 162 353
rect 172 352 192 493
rect 171 351 192 352
rect 134 349 163 351
rect 170 350 192 351
rect 169 349 192 350
rect 135 347 164 349
rect 168 348 192 349
rect 167 347 192 348
rect 136 346 165 347
rect 166 346 192 347
rect 136 345 192 346
rect 137 343 192 345
rect 138 341 192 343
rect 139 339 192 341
rect 140 337 192 339
rect 141 335 192 337
rect 142 333 192 335
rect 212 352 232 493
rect 272 492 492 493
rect 271 491 492 492
rect 270 490 492 491
rect 269 489 492 490
rect 268 488 492 489
rect 267 487 492 488
rect 266 486 492 487
rect 265 485 492 486
rect 264 484 492 485
rect 263 483 492 484
rect 262 482 492 483
rect 261 481 492 482
rect 260 480 492 481
rect 259 479 492 480
rect 258 478 492 479
rect 257 477 492 478
rect 256 476 492 477
rect 255 475 492 476
rect 254 474 492 475
rect 253 473 492 474
rect 252 472 291 473
rect 252 471 290 472
rect 252 470 289 471
rect 252 469 288 470
rect 252 468 287 469
rect 252 467 286 468
rect 252 466 285 467
rect 252 465 284 466
rect 252 464 283 465
rect 252 463 282 464
rect 252 462 281 463
rect 252 461 280 462
rect 252 460 279 461
rect 252 459 278 460
rect 252 458 277 459
rect 252 457 276 458
rect 252 456 275 457
rect 252 455 274 456
rect 252 454 273 455
rect 252 432 272 454
rect 252 431 273 432
rect 252 430 274 431
rect 252 429 275 430
rect 252 428 276 429
rect 252 427 277 428
rect 252 426 278 427
rect 252 425 279 426
rect 252 424 280 425
rect 252 423 281 424
rect 252 422 282 423
rect 252 421 283 422
rect 252 420 284 421
rect 252 419 285 420
rect 252 418 286 419
rect 252 417 287 418
rect 252 416 288 417
rect 252 415 289 416
rect 252 414 290 415
rect 252 413 291 414
rect 253 412 372 413
rect 254 411 373 412
rect 255 410 374 411
rect 256 409 375 410
rect 257 408 376 409
rect 258 407 377 408
rect 259 406 378 407
rect 260 405 379 406
rect 261 404 380 405
rect 262 403 381 404
rect 263 402 382 403
rect 264 401 383 402
rect 265 400 384 401
rect 266 399 385 400
rect 267 398 386 399
rect 268 397 387 398
rect 269 396 388 397
rect 270 395 389 396
rect 271 394 390 395
rect 272 393 391 394
rect 353 392 392 393
rect 354 391 392 392
rect 355 390 392 391
rect 356 389 392 390
rect 357 388 392 389
rect 358 387 392 388
rect 359 386 392 387
rect 360 385 392 386
rect 361 384 392 385
rect 362 383 392 384
rect 363 382 392 383
rect 364 381 392 382
rect 365 380 392 381
rect 366 379 392 380
rect 367 378 392 379
rect 368 377 392 378
rect 369 376 392 377
rect 370 375 392 376
rect 371 374 392 375
rect 372 352 392 374
rect 212 351 233 352
rect 371 351 392 352
rect 212 350 234 351
rect 370 350 392 351
rect 212 349 235 350
rect 369 349 392 350
rect 212 348 236 349
rect 368 348 392 349
rect 212 347 237 348
rect 367 347 392 348
rect 212 346 238 347
rect 366 346 392 347
rect 212 345 239 346
rect 365 345 392 346
rect 212 344 240 345
rect 364 344 392 345
rect 212 343 241 344
rect 363 343 392 344
rect 212 342 242 343
rect 362 342 392 343
rect 212 341 243 342
rect 361 341 392 342
rect 212 340 244 341
rect 360 340 392 341
rect 212 339 245 340
rect 359 339 392 340
rect 212 338 246 339
rect 358 338 392 339
rect 212 337 247 338
rect 357 337 392 338
rect 212 336 248 337
rect 356 336 392 337
rect 212 335 249 336
rect 355 335 392 336
rect 212 334 250 335
rect 354 334 392 335
rect 212 333 251 334
rect 353 333 392 334
rect 143 332 191 333
rect 213 332 392 333
rect 143 331 190 332
rect 214 331 390 332
rect 144 330 189 331
rect 215 330 389 331
rect 144 329 188 330
rect 216 329 388 330
rect 145 328 187 329
rect 217 328 387 329
rect 145 327 186 328
rect 218 327 386 328
rect 146 326 185 327
rect 219 326 385 327
rect 146 325 184 326
rect 220 325 384 326
rect 147 324 183 325
rect 221 324 383 325
rect 147 323 182 324
rect 222 323 382 324
rect 148 322 181 323
rect 223 322 381 323
rect 148 321 180 322
rect 224 321 380 322
rect 149 320 179 321
rect 225 320 379 321
rect 149 319 178 320
rect 226 319 378 320
rect 150 318 177 319
rect 227 318 377 319
rect 150 317 176 318
rect 228 317 376 318
rect 151 316 175 317
rect 229 316 375 317
rect 151 315 174 316
rect 230 315 374 316
rect 152 314 173 315
rect 231 314 373 315
rect 152 313 172 314
rect 232 313 372 314
rect 412 313 432 473
rect 508 419 658 449
rect 868 419 988 449
rect 568 329 598 419
rect 688 418 718 419
rect 808 418 838 419
rect 688 417 719 418
rect 807 417 838 418
rect 688 416 720 417
rect 806 416 838 417
rect 688 415 721 416
rect 805 415 838 416
rect 688 414 722 415
rect 804 414 838 415
rect 688 413 723 414
rect 803 413 838 414
rect 688 412 724 413
rect 802 412 838 413
rect 688 411 725 412
rect 801 411 838 412
rect 688 410 726 411
rect 800 410 838 411
rect 688 409 727 410
rect 799 409 838 410
rect 688 408 728 409
rect 798 408 838 409
rect 688 407 729 408
rect 797 407 838 408
rect 688 406 730 407
rect 796 406 838 407
rect 688 405 731 406
rect 795 405 838 406
rect 688 404 732 405
rect 794 404 838 405
rect 688 403 733 404
rect 793 403 838 404
rect 688 402 734 403
rect 792 402 838 403
rect 688 401 735 402
rect 791 401 838 402
rect 688 400 736 401
rect 790 400 838 401
rect 688 399 737 400
rect 789 399 838 400
rect 688 398 738 399
rect 788 398 838 399
rect 688 397 739 398
rect 787 397 838 398
rect 688 396 740 397
rect 786 396 838 397
rect 688 395 741 396
rect 785 395 838 396
rect 688 394 742 395
rect 784 394 838 395
rect 688 393 743 394
rect 783 393 838 394
rect 688 392 744 393
rect 782 392 838 393
rect 688 391 745 392
rect 781 391 838 392
rect 688 390 746 391
rect 780 390 838 391
rect 688 389 747 390
rect 779 389 838 390
rect 688 388 748 389
rect 778 388 838 389
rect 688 387 749 388
rect 777 387 838 388
rect 688 386 750 387
rect 776 386 838 387
rect 688 385 751 386
rect 775 385 838 386
rect 688 384 752 385
rect 774 384 838 385
rect 688 383 753 384
rect 773 383 838 384
rect 688 382 754 383
rect 772 382 838 383
rect 688 381 755 382
rect 771 381 838 382
rect 688 380 756 381
rect 770 380 838 381
rect 688 379 757 380
rect 769 379 838 380
rect 688 378 758 379
rect 768 378 838 379
rect 688 377 759 378
rect 767 377 838 378
rect 688 376 760 377
rect 766 376 838 377
rect 688 375 761 376
rect 765 375 838 376
rect 688 374 762 375
rect 764 374 838 375
rect 688 359 838 374
rect 868 389 898 419
rect 868 359 988 389
rect 508 299 658 329
rect 503 284 518 289
rect 520 286 525 289
rect 508 274 513 284
rect 520 283 527 286
rect 520 280 529 283
rect 530 280 535 289
rect 537 284 552 289
rect 554 284 569 289
rect 571 284 586 289
rect 588 284 603 289
rect 520 278 535 280
rect 503 269 518 274
rect 520 269 525 278
rect 526 275 535 278
rect 528 272 535 275
rect 530 269 535 272
rect 542 269 547 284
rect 554 281 559 284
rect 554 276 564 281
rect 554 274 559 276
rect 571 274 576 284
rect 588 281 593 284
rect 598 281 603 284
rect 579 276 586 281
rect 581 274 586 276
rect 554 269 569 274
rect 571 269 586 274
rect 588 276 603 281
rect 605 284 620 289
rect 622 284 637 289
rect 639 284 654 289
rect 658 288 668 289
rect 658 287 670 288
rect 658 284 672 287
rect 605 281 610 284
rect 615 281 620 284
rect 605 276 620 281
rect 588 275 601 276
rect 588 274 602 275
rect 588 269 593 274
rect 594 273 603 274
rect 595 272 603 273
rect 596 271 603 272
rect 597 270 603 271
rect 598 269 603 270
rect 605 269 610 276
rect 615 269 620 276
rect 627 269 632 284
rect 639 281 644 284
rect 639 276 649 281
rect 639 274 644 276
rect 658 274 663 284
rect 665 283 673 284
rect 667 282 673 283
rect 668 276 673 282
rect 667 275 673 276
rect 665 274 673 275
rect 639 269 654 274
rect 658 271 672 274
rect 658 270 670 271
rect 658 269 668 270
rect 688 269 718 359
rect 719 358 807 359
rect 720 357 806 358
rect 721 356 805 357
rect 722 355 804 356
rect 723 354 803 355
rect 724 353 802 354
rect 725 352 801 353
rect 726 351 800 352
rect 727 350 799 351
rect 728 349 798 350
rect 729 348 797 349
rect 730 347 796 348
rect 731 346 795 347
rect 732 345 794 346
rect 733 344 793 345
rect 734 343 792 344
rect 735 342 791 343
rect 736 341 790 342
rect 737 340 789 341
rect 738 339 788 340
rect 739 338 787 339
rect 740 337 786 338
rect 741 336 785 337
rect 742 335 784 336
rect 743 334 783 335
rect 744 333 782 334
rect 745 332 781 333
rect 746 331 780 332
rect 747 330 779 331
rect 748 329 778 330
rect 749 328 777 329
rect 750 327 776 328
rect 751 326 775 327
rect 752 325 774 326
rect 753 324 773 325
rect 754 323 772 324
rect 755 322 771 323
rect 756 321 770 322
rect 757 320 769 321
rect 758 319 768 320
rect 759 318 767 319
rect 760 317 766 318
rect 761 316 765 317
rect 762 315 764 316
rect 808 269 838 359
rect 958 329 988 359
rect 868 299 988 329
rect 863 284 878 289
rect 880 286 885 289
rect 895 286 900 289
rect 880 284 887 286
rect 863 281 868 284
rect 882 283 887 284
rect 893 284 900 286
rect 902 284 917 289
rect 919 284 934 289
rect 936 284 951 289
rect 953 286 958 289
rect 968 286 973 289
rect 893 283 898 284
rect 882 281 889 283
rect 863 276 878 281
rect 884 280 889 281
rect 891 281 898 283
rect 902 281 907 284
rect 891 280 896 281
rect 884 278 896 280
rect 873 274 878 276
rect 886 275 894 278
rect 902 276 917 281
rect 863 269 878 274
rect 888 269 893 275
rect 912 274 917 276
rect 902 269 917 274
rect 924 269 929 284
rect 936 281 941 284
rect 953 283 960 286
rect 966 283 973 286
rect 936 276 946 281
rect 953 280 962 283
rect 964 280 973 283
rect 953 278 973 280
rect 936 274 941 276
rect 936 269 951 274
rect 953 269 958 278
rect 959 275 967 278
rect 968 269 973 278
rect 975 284 990 289
rect 975 281 980 284
rect 975 276 990 281
rect 985 274 990 276
rect 975 269 990 274
rect 666 251 671 254
rect 681 251 686 254
rect 666 248 673 251
rect 679 248 686 251
rect 666 245 675 248
rect 677 245 686 248
rect 666 243 686 245
rect 666 234 671 243
rect 672 240 680 243
rect 681 234 686 243
rect 688 249 703 254
rect 705 249 720 254
rect 688 246 693 249
rect 705 246 710 249
rect 715 246 720 249
rect 688 241 698 246
rect 705 241 720 246
rect 722 249 737 254
rect 722 246 727 249
rect 722 241 737 246
rect 688 239 693 241
rect 688 234 703 239
rect 705 234 710 241
rect 715 234 720 241
rect 732 239 737 241
rect 722 234 737 239
rect 739 239 744 254
rect 749 239 754 254
rect 739 234 754 239
rect 756 249 771 254
rect 756 246 761 249
rect 766 246 771 249
rect 756 241 771 246
rect 774 249 789 254
rect 791 251 796 254
rect 806 251 811 254
rect 774 246 779 249
rect 791 248 798 251
rect 804 248 811 251
rect 774 241 784 246
rect 791 245 800 248
rect 802 245 811 248
rect 791 243 811 245
rect 756 240 769 241
rect 756 239 770 240
rect 774 239 779 241
rect 756 234 761 239
rect 762 238 771 239
rect 763 237 771 238
rect 764 236 771 237
rect 765 235 771 236
rect 766 234 771 235
rect 774 234 789 239
rect 791 234 796 243
rect 797 240 805 243
rect 806 234 811 243
rect 813 249 828 254
rect 830 251 835 254
rect 813 246 818 249
rect 830 248 837 251
rect 813 241 823 246
rect 830 245 839 248
rect 840 245 845 254
rect 847 249 862 254
rect 830 243 845 245
rect 813 239 818 241
rect 813 234 828 239
rect 830 234 835 243
rect 836 240 845 243
rect 838 237 845 240
rect 840 234 845 237
rect 852 234 857 249
<< metal1 >>
rect 105 210 155 220
rect 105 170 115 210
rect 125 170 135 210
rect 145 170 155 210
rect 165 210 195 220
rect 205 210 255 220
rect 165 200 175 210
rect 165 190 185 200
rect 165 180 175 190
rect 165 170 195 180
rect 205 170 215 210
rect 225 170 235 210
rect 245 170 255 210
rect 265 210 295 220
rect 265 200 275 210
rect 265 190 295 200
rect 285 180 295 190
rect 265 170 295 180
rect 345 180 355 220
rect 385 210 415 220
rect 425 210 455 220
rect 395 180 405 210
rect 425 200 435 210
rect 445 200 455 210
rect 425 190 455 200
rect 425 180 435 190
rect 445 180 455 190
rect 345 170 375 180
rect 385 170 415 180
rect 425 170 455 180
rect 465 215 490 220
rect 465 210 495 215
rect 465 200 475 210
rect 485 200 495 210
rect 505 210 535 220
rect 505 200 515 210
rect 525 200 535 210
rect 465 190 490 200
rect 505 190 535 200
rect 465 170 475 190
rect 485 170 495 190
rect 505 170 515 190
rect 525 170 535 190
rect 545 215 570 220
rect 545 210 575 215
rect 545 200 555 210
rect 565 200 575 210
rect 585 200 595 220
rect 605 200 615 220
rect 545 190 570 200
rect 585 190 615 200
rect 545 170 555 190
rect 565 170 575 190
rect 595 170 605 190
use open-80x80 2_0
timestamp 760840415
transform 1 0 -210 0 1 259
box 488 -239 568 -159
use open-oxide-80x80 3_0
timestamp 760840453
transform 1 0 -359 0 1 142
box 637 -242 717 -162
use thermal-converter 4_0
timestamp 760840748
transform 1 0 461 0 1 10
box -16 -110 134 110
use thermal-actuator 5_0
timestamp 760840666
transform 1 0 675 0 1 -100
box 0 0 90 220
use pixel-80x80 6_0
timestamp 760840526
transform 1 0 -430 0 1 -336
box 497 -3 587 87
use pixel-160x160 7_0
timestamp 760840608
transform 1 0 -80 0 1 -367
box 288 -12 458 158
use micro-hot-plate 8_0
timestamp 760840982
transform 1 0 420 0 1 -430
box 0 0 260 266
use gas-sensor 9_0
timestamp 760840948
transform 1 0 720 0 1 -430
box 0 0 260 266
<< end >>
