magic
tech scmos
timestamp 500618087
<< error_s >>
rect 49 6 50 8
<< polysilicon >>
rect 19 15 21 46
rect 28 15 30 46
rect 33 15 35 46
rect 21 -37 23 -6
rect 25 -37 27 -6
rect 33 -37 35 -6
<< ndiffusion >>
rect 15 15 17 46
<< metal1 >>
rect 50 10 64 13
rect -6 1 3 4
rect -6 -6 3 -2
rect 50 -6 65 -2
use tut3e tut3e_0
timestamp 500618087
transform 1 0 3 0 1 -6
box 0 0 47 21
<< labels >>
rlabel space 72 4 72 4 7 Point here
<< end >>
