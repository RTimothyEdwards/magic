magic
tech scmos
timestamp 760840415
<< substrateopen >>
rect 488 -239 568 -159
<< end >>
