magic
tech scmos
timestamp 760840948
<< polysilicon >>
rect 250 265 260 266
rect 249 264 260 265
rect 248 263 260 264
rect 247 262 253 263
rect 246 261 253 262
rect 245 260 253 261
rect 244 259 253 260
rect 257 259 260 263
rect 243 258 260 259
rect 242 257 260 258
rect 241 256 260 257
rect 240 255 259 256
rect 239 254 258 255
rect 238 253 257 254
rect 237 252 256 253
rect 236 251 255 252
rect 235 250 254 251
rect 234 249 253 250
rect 233 248 252 249
rect 232 247 251 248
rect 231 246 250 247
rect 230 245 249 246
rect 229 244 248 245
rect 228 243 247 244
rect 227 242 246 243
rect 226 241 245 242
rect 225 240 244 241
rect 224 239 243 240
rect 223 238 242 239
rect 222 237 241 238
rect 221 236 240 237
rect 220 235 239 236
rect 219 234 238 235
rect 218 233 237 234
rect 217 232 236 233
rect 216 231 235 232
rect 215 230 234 231
rect 214 229 233 230
rect 213 228 232 229
rect 212 227 231 228
rect 211 226 230 227
rect 210 225 229 226
rect 209 224 228 225
rect 208 223 227 224
rect 207 222 226 223
rect 206 221 225 222
rect 205 220 224 221
rect 204 219 223 220
rect 203 218 222 219
rect 202 217 221 218
rect 201 216 220 217
rect 200 215 219 216
rect 199 214 218 215
rect 198 213 217 214
rect 197 212 216 213
rect 196 211 215 212
rect 195 210 214 211
rect 194 209 213 210
rect 193 208 212 209
rect 192 207 211 208
rect 191 206 210 207
rect 190 205 209 206
rect 189 204 208 205
rect 188 203 207 204
rect 187 202 206 203
rect 186 201 205 202
rect 185 200 204 201
rect 184 199 203 200
rect 183 198 202 199
rect 182 197 201 198
rect 181 196 200 197
rect 180 195 199 196
rect 179 194 198 195
rect 178 193 197 194
rect 177 192 196 193
rect 176 191 195 192
rect 175 190 194 191
rect 174 189 193 190
rect 173 188 192 189
rect 172 187 191 188
rect 171 186 190 187
rect 170 185 189 186
rect 169 184 188 185
rect 168 183 187 184
rect 167 182 186 183
rect 166 181 185 182
rect 165 180 184 181
rect 164 179 183 180
rect 163 178 182 179
rect 162 177 181 178
rect 162 176 180 177
rect 90 175 179 176
rect 90 174 178 175
rect 90 173 177 174
rect 90 172 176 173
rect 90 171 175 172
rect 90 170 174 171
rect 90 169 173 170
rect 90 168 172 169
rect 90 164 98 168
rect 90 156 170 164
rect 162 152 170 156
rect 90 144 170 152
rect 90 140 98 144
rect 90 132 170 140
rect 162 128 170 132
rect 90 120 170 128
rect 90 116 98 120
rect 90 108 170 116
rect 162 104 170 108
rect 88 103 170 104
rect 87 102 170 103
rect 86 101 170 102
rect 85 100 170 101
rect 84 99 170 100
rect 83 98 170 99
rect 82 97 170 98
rect 81 96 170 97
rect 80 95 98 96
rect 79 94 98 95
rect 78 93 97 94
rect 77 92 96 93
rect 76 91 95 92
rect 75 90 94 91
rect 74 89 93 90
rect 73 88 92 89
rect 72 87 91 88
rect 71 86 90 87
rect 70 85 89 86
rect 69 84 88 85
rect 68 83 87 84
rect 67 82 86 83
rect 66 81 85 82
rect 65 80 84 81
rect 64 79 83 80
rect 63 78 82 79
rect 62 77 81 78
rect 61 76 80 77
rect 60 75 79 76
rect 59 74 78 75
rect 58 73 77 74
rect 57 72 76 73
rect 56 71 75 72
rect 55 70 74 71
rect 54 69 73 70
rect 53 68 72 69
rect 52 67 71 68
rect 51 66 70 67
rect 50 65 69 66
rect 49 64 68 65
rect 48 63 67 64
rect 47 62 66 63
rect 46 61 65 62
rect 45 60 64 61
rect 44 59 63 60
rect 43 58 62 59
rect 42 57 61 58
rect 41 56 60 57
rect 40 55 59 56
rect 39 54 58 55
rect 38 53 57 54
rect 37 52 56 53
rect 36 51 55 52
rect 35 50 54 51
rect 34 49 53 50
rect 33 48 52 49
rect 32 47 51 48
rect 31 46 50 47
rect 30 45 49 46
rect 29 44 48 45
rect 28 43 47 44
rect 27 42 46 43
rect 26 41 45 42
rect 25 40 44 41
rect 24 39 43 40
rect 23 38 42 39
rect 22 37 41 38
rect 21 36 40 37
rect 20 35 39 36
rect 19 34 38 35
rect 18 33 37 34
rect 17 32 36 33
rect 16 31 35 32
rect 15 30 34 31
rect 14 29 33 30
rect 13 28 32 29
rect 12 27 31 28
rect 11 26 30 27
rect 10 25 29 26
rect 9 24 28 25
rect 8 23 27 24
rect 7 22 26 23
rect 6 21 25 22
rect 5 20 24 21
rect 4 19 23 20
rect 3 18 22 19
rect 2 17 21 18
rect 1 16 20 17
rect 0 15 19 16
rect 0 14 18 15
rect 0 13 17 14
rect 0 9 3 13
rect 7 12 16 13
rect 7 11 15 12
rect 7 10 14 11
rect 7 9 13 10
rect 0 8 12 9
rect 0 7 11 8
rect 0 6 10 7
<< metal1 >>
rect 250 263 260 266
rect 250 259 253 263
rect 257 259 260 263
rect 250 256 260 259
rect 0 240 30 246
rect 230 240 260 246
rect 0 239 31 240
rect 229 239 260 240
rect 0 238 32 239
rect 228 238 260 239
rect 0 237 33 238
rect 227 237 260 238
rect 0 236 34 237
rect 226 236 260 237
rect 26 235 35 236
rect 225 235 234 236
rect 27 234 36 235
rect 224 234 233 235
rect 28 233 37 234
rect 223 233 232 234
rect 29 232 38 233
rect 222 232 231 233
rect 30 231 39 232
rect 221 231 230 232
rect 31 230 40 231
rect 220 230 229 231
rect 32 229 41 230
rect 219 229 228 230
rect 33 228 42 229
rect 218 228 227 229
rect 34 227 43 228
rect 217 227 226 228
rect 35 226 44 227
rect 216 226 225 227
rect 36 225 45 226
rect 215 225 224 226
rect 37 224 46 225
rect 214 224 223 225
rect 38 223 47 224
rect 213 223 222 224
rect 39 222 48 223
rect 212 222 221 223
rect 40 221 49 222
rect 211 221 220 222
rect 41 220 50 221
rect 210 220 219 221
rect 42 219 51 220
rect 209 219 218 220
rect 43 218 52 219
rect 208 218 217 219
rect 44 217 53 218
rect 207 217 216 218
rect 45 216 54 217
rect 206 216 215 217
rect 46 215 55 216
rect 205 215 214 216
rect 47 214 56 215
rect 204 214 213 215
rect 48 213 57 214
rect 203 213 212 214
rect 49 212 58 213
rect 202 212 211 213
rect 50 211 59 212
rect 201 211 210 212
rect 51 210 60 211
rect 200 210 209 211
rect 52 209 61 210
rect 199 209 208 210
rect 53 208 62 209
rect 198 208 207 209
rect 54 207 63 208
rect 197 207 206 208
rect 55 206 64 207
rect 196 206 205 207
rect 56 205 65 206
rect 195 205 204 206
rect 57 204 66 205
rect 194 204 203 205
rect 58 203 67 204
rect 193 203 202 204
rect 59 202 68 203
rect 192 202 201 203
rect 60 201 69 202
rect 191 201 200 202
rect 61 200 70 201
rect 190 200 199 201
rect 62 199 71 200
rect 189 199 198 200
rect 63 198 72 199
rect 188 198 197 199
rect 64 197 73 198
rect 187 197 196 198
rect 65 196 74 197
rect 186 196 195 197
rect 66 195 75 196
rect 185 195 194 196
rect 67 194 76 195
rect 184 194 193 195
rect 68 193 77 194
rect 183 193 192 194
rect 69 192 78 193
rect 182 192 191 193
rect 70 191 79 192
rect 181 191 190 192
rect 71 190 80 191
rect 180 190 189 191
rect 72 189 81 190
rect 179 189 188 190
rect 73 188 82 189
rect 178 188 187 189
rect 74 187 83 188
rect 177 187 186 188
rect 75 186 84 187
rect 176 186 185 187
rect 76 185 85 186
rect 175 185 184 186
rect 77 184 86 185
rect 174 184 183 185
rect 78 183 87 184
rect 173 183 182 184
rect 79 182 88 183
rect 172 182 181 183
rect 80 181 89 182
rect 171 181 180 182
rect 81 180 179 181
rect 82 179 178 180
rect 83 178 177 179
rect 84 177 176 178
rect 85 95 175 177
rect 84 94 176 95
rect 83 93 177 94
rect 82 92 178 93
rect 81 91 179 92
rect 80 90 89 91
rect 171 90 180 91
rect 79 89 88 90
rect 172 89 181 90
rect 78 88 87 89
rect 173 88 182 89
rect 77 87 86 88
rect 174 87 183 88
rect 76 86 85 87
rect 175 86 184 87
rect 75 85 84 86
rect 176 85 185 86
rect 74 84 83 85
rect 177 84 186 85
rect 73 83 82 84
rect 178 83 187 84
rect 72 82 81 83
rect 179 82 188 83
rect 71 81 80 82
rect 180 81 189 82
rect 70 80 79 81
rect 181 80 190 81
rect 69 79 78 80
rect 182 79 191 80
rect 68 78 77 79
rect 183 78 192 79
rect 67 77 76 78
rect 184 77 193 78
rect 66 76 75 77
rect 185 76 194 77
rect 65 75 74 76
rect 186 75 195 76
rect 64 74 73 75
rect 187 74 196 75
rect 63 73 72 74
rect 188 73 197 74
rect 62 72 71 73
rect 189 72 198 73
rect 61 71 70 72
rect 190 71 199 72
rect 60 70 69 71
rect 191 70 200 71
rect 59 69 68 70
rect 192 69 201 70
rect 58 68 67 69
rect 193 68 202 69
rect 57 67 66 68
rect 194 67 203 68
rect 56 66 65 67
rect 195 66 204 67
rect 55 65 64 66
rect 196 65 205 66
rect 54 64 63 65
rect 197 64 206 65
rect 53 63 62 64
rect 198 63 207 64
rect 52 62 61 63
rect 199 62 208 63
rect 51 61 60 62
rect 200 61 209 62
rect 50 60 59 61
rect 201 60 210 61
rect 49 59 58 60
rect 202 59 211 60
rect 48 58 57 59
rect 203 58 212 59
rect 47 57 56 58
rect 204 57 213 58
rect 46 56 55 57
rect 205 56 214 57
rect 45 55 54 56
rect 206 55 215 56
rect 44 54 53 55
rect 207 54 216 55
rect 43 53 52 54
rect 208 53 217 54
rect 42 52 51 53
rect 209 52 218 53
rect 41 51 50 52
rect 210 51 219 52
rect 40 50 49 51
rect 211 50 220 51
rect 39 49 48 50
rect 212 49 221 50
rect 38 48 47 49
rect 213 48 222 49
rect 37 47 46 48
rect 214 47 223 48
rect 36 46 45 47
rect 215 46 224 47
rect 35 45 44 46
rect 216 45 225 46
rect 34 44 43 45
rect 217 44 226 45
rect 33 43 42 44
rect 218 43 227 44
rect 32 42 41 43
rect 219 42 228 43
rect 31 41 40 42
rect 220 41 229 42
rect 30 40 39 41
rect 221 40 230 41
rect 29 39 38 40
rect 222 39 231 40
rect 28 38 37 39
rect 223 38 232 39
rect 27 37 36 38
rect 224 37 233 38
rect 26 36 35 37
rect 225 36 234 37
rect 0 35 34 36
rect 226 35 260 36
rect 0 34 33 35
rect 227 34 260 35
rect 0 33 32 34
rect 228 33 260 34
rect 0 32 31 33
rect 229 32 260 33
rect 0 26 30 32
rect 230 26 260 32
rect 0 13 10 16
rect 0 9 3 13
rect 7 9 10 13
rect 0 0 10 9
<< metal2 >>
rect 20 240 30 266
rect 230 240 240 266
rect 20 239 31 240
rect 229 239 240 240
rect 20 238 32 239
rect 228 238 240 239
rect 20 237 33 238
rect 227 237 240 238
rect 20 236 34 237
rect 226 236 240 237
rect 26 235 35 236
rect 225 235 234 236
rect 27 234 36 235
rect 224 234 233 235
rect 28 233 37 234
rect 223 233 232 234
rect 29 232 38 233
rect 222 232 231 233
rect 30 231 39 232
rect 221 231 230 232
rect 31 230 40 231
rect 220 230 229 231
rect 32 229 41 230
rect 219 229 228 230
rect 33 228 42 229
rect 218 228 227 229
rect 34 227 43 228
rect 217 227 226 228
rect 35 226 44 227
rect 216 226 225 227
rect 36 225 45 226
rect 215 225 224 226
rect 37 224 46 225
rect 214 224 223 225
rect 38 223 47 224
rect 213 223 222 224
rect 39 222 48 223
rect 212 222 221 223
rect 40 221 49 222
rect 211 221 220 222
rect 41 220 50 221
rect 210 220 219 221
rect 42 219 51 220
rect 209 219 218 220
rect 43 218 52 219
rect 208 218 217 219
rect 44 217 53 218
rect 207 217 216 218
rect 45 216 54 217
rect 206 216 215 217
rect 46 215 55 216
rect 205 215 214 216
rect 47 214 56 215
rect 204 214 213 215
rect 48 213 57 214
rect 203 213 212 214
rect 49 212 58 213
rect 202 212 211 213
rect 50 211 59 212
rect 201 211 210 212
rect 51 210 60 211
rect 200 210 209 211
rect 52 209 61 210
rect 199 209 208 210
rect 53 208 62 209
rect 198 208 207 209
rect 54 207 63 208
rect 197 207 206 208
rect 55 206 64 207
rect 196 206 205 207
rect 56 205 65 206
rect 195 205 204 206
rect 57 204 66 205
rect 194 204 203 205
rect 58 203 67 204
rect 193 203 202 204
rect 59 202 68 203
rect 192 202 201 203
rect 60 201 69 202
rect 191 201 200 202
rect 61 200 70 201
rect 190 200 199 201
rect 62 199 71 200
rect 189 199 198 200
rect 63 198 72 199
rect 188 198 197 199
rect 64 197 73 198
rect 187 197 196 198
rect 65 196 74 197
rect 186 196 195 197
rect 66 195 75 196
rect 185 195 194 196
rect 67 194 76 195
rect 184 194 193 195
rect 68 193 77 194
rect 183 193 192 194
rect 69 192 78 193
rect 182 192 191 193
rect 70 191 79 192
rect 181 191 190 192
rect 71 190 80 191
rect 180 190 189 191
rect 72 189 81 190
rect 179 189 188 190
rect 73 188 82 189
rect 178 188 187 189
rect 74 187 83 188
rect 177 187 186 188
rect 75 186 84 187
rect 176 186 185 187
rect 76 185 85 186
rect 175 185 184 186
rect 77 184 86 185
rect 174 184 183 185
rect 78 183 87 184
rect 173 183 182 184
rect 79 182 88 183
rect 172 182 181 183
rect 80 181 89 182
rect 171 181 180 182
rect 81 180 90 181
rect 170 180 179 181
rect 82 179 91 180
rect 169 179 178 180
rect 83 178 92 179
rect 168 178 177 179
rect 84 177 93 178
rect 167 177 176 178
rect 85 176 94 177
rect 166 176 175 177
rect 86 175 125 176
rect 87 174 125 175
rect 88 173 125 174
rect 89 172 125 173
rect 90 141 125 172
rect 135 175 174 176
rect 135 174 173 175
rect 135 173 172 174
rect 135 172 171 173
rect 135 141 170 172
rect 90 100 125 131
rect 89 99 125 100
rect 88 98 125 99
rect 87 97 125 98
rect 86 96 125 97
rect 135 100 170 131
rect 135 99 171 100
rect 135 98 172 99
rect 135 97 173 98
rect 135 96 174 97
rect 85 95 94 96
rect 166 95 175 96
rect 84 94 93 95
rect 167 94 176 95
rect 83 93 92 94
rect 168 93 177 94
rect 82 92 91 93
rect 169 92 178 93
rect 81 91 90 92
rect 170 91 179 92
rect 80 90 89 91
rect 171 90 180 91
rect 79 89 88 90
rect 172 89 181 90
rect 78 88 87 89
rect 173 88 182 89
rect 77 87 86 88
rect 174 87 183 88
rect 76 86 85 87
rect 175 86 184 87
rect 75 85 84 86
rect 176 85 185 86
rect 74 84 83 85
rect 177 84 186 85
rect 73 83 82 84
rect 178 83 187 84
rect 72 82 81 83
rect 179 82 188 83
rect 71 81 80 82
rect 180 81 189 82
rect 70 80 79 81
rect 181 80 190 81
rect 69 79 78 80
rect 182 79 191 80
rect 68 78 77 79
rect 183 78 192 79
rect 67 77 76 78
rect 184 77 193 78
rect 66 76 75 77
rect 185 76 194 77
rect 65 75 74 76
rect 186 75 195 76
rect 64 74 73 75
rect 187 74 196 75
rect 63 73 72 74
rect 188 73 197 74
rect 62 72 71 73
rect 189 72 198 73
rect 61 71 70 72
rect 190 71 199 72
rect 60 70 69 71
rect 191 70 200 71
rect 59 69 68 70
rect 192 69 201 70
rect 58 68 67 69
rect 193 68 202 69
rect 57 67 66 68
rect 194 67 203 68
rect 56 66 65 67
rect 195 66 204 67
rect 55 65 64 66
rect 196 65 205 66
rect 54 64 63 65
rect 197 64 206 65
rect 53 63 62 64
rect 198 63 207 64
rect 52 62 61 63
rect 199 62 208 63
rect 51 61 60 62
rect 200 61 209 62
rect 50 60 59 61
rect 201 60 210 61
rect 49 59 58 60
rect 202 59 211 60
rect 48 58 57 59
rect 203 58 212 59
rect 47 57 56 58
rect 204 57 213 58
rect 46 56 55 57
rect 205 56 214 57
rect 45 55 54 56
rect 206 55 215 56
rect 44 54 53 55
rect 207 54 216 55
rect 43 53 52 54
rect 208 53 217 54
rect 42 52 51 53
rect 209 52 218 53
rect 41 51 50 52
rect 210 51 219 52
rect 40 50 49 51
rect 211 50 220 51
rect 39 49 48 50
rect 212 49 221 50
rect 38 48 47 49
rect 213 48 222 49
rect 37 47 46 48
rect 214 47 223 48
rect 36 46 45 47
rect 215 46 224 47
rect 35 45 44 46
rect 216 45 225 46
rect 34 44 43 45
rect 217 44 226 45
rect 33 43 42 44
rect 218 43 227 44
rect 32 42 41 43
rect 219 42 228 43
rect 31 41 40 42
rect 220 41 229 42
rect 30 40 39 41
rect 221 40 230 41
rect 29 39 38 40
rect 222 39 231 40
rect 28 38 37 39
rect 223 38 232 39
rect 27 37 36 38
rect 224 37 233 38
rect 26 36 35 37
rect 225 36 234 37
rect 20 35 34 36
rect 226 35 240 36
rect 20 34 33 35
rect 227 34 240 35
rect 20 33 32 34
rect 228 33 240 34
rect 20 32 31 33
rect 229 32 240 33
rect 20 6 30 32
rect 230 6 240 32
<< polycontact >>
rect 253 259 257 263
rect 3 9 7 13
<< substrateopen >>
rect 50 235 210 236
rect 51 234 209 235
rect 52 233 208 234
rect 53 232 207 233
rect 54 231 206 232
rect 55 230 205 231
rect 56 229 204 230
rect 57 228 203 229
rect 58 227 202 228
rect 59 226 201 227
rect 60 225 200 226
rect 61 224 199 225
rect 62 223 198 224
rect 63 222 197 223
rect 64 221 196 222
rect 65 220 195 221
rect 66 219 194 220
rect 67 218 193 219
rect 68 217 192 218
rect 69 216 191 217
rect 30 215 31 216
rect 70 215 190 216
rect 229 215 230 216
rect 30 214 32 215
rect 71 214 189 215
rect 228 214 230 215
rect 30 213 33 214
rect 72 213 188 214
rect 227 213 230 214
rect 30 212 34 213
rect 73 212 187 213
rect 226 212 230 213
rect 30 211 35 212
rect 74 211 186 212
rect 225 211 230 212
rect 30 210 36 211
rect 75 210 185 211
rect 224 210 230 211
rect 30 209 37 210
rect 76 209 184 210
rect 223 209 230 210
rect 30 208 38 209
rect 77 208 183 209
rect 222 208 230 209
rect 30 207 39 208
rect 78 207 182 208
rect 221 207 230 208
rect 30 206 40 207
rect 79 206 181 207
rect 220 206 230 207
rect 30 205 41 206
rect 80 205 180 206
rect 219 205 230 206
rect 30 204 42 205
rect 81 204 179 205
rect 218 204 230 205
rect 30 203 43 204
rect 82 203 178 204
rect 217 203 230 204
rect 30 202 44 203
rect 83 202 177 203
rect 216 202 230 203
rect 30 201 45 202
rect 84 201 176 202
rect 215 201 230 202
rect 30 200 46 201
rect 85 200 175 201
rect 214 200 230 201
rect 30 199 47 200
rect 86 199 174 200
rect 213 199 230 200
rect 30 198 48 199
rect 87 198 173 199
rect 212 198 230 199
rect 30 197 49 198
rect 88 197 172 198
rect 211 197 230 198
rect 30 196 50 197
rect 89 196 171 197
rect 210 196 230 197
rect 30 195 51 196
rect 90 195 170 196
rect 209 195 230 196
rect 30 194 52 195
rect 91 194 169 195
rect 208 194 230 195
rect 30 193 53 194
rect 92 193 168 194
rect 207 193 230 194
rect 30 192 54 193
rect 93 192 167 193
rect 206 192 230 193
rect 30 191 55 192
rect 94 191 166 192
rect 205 191 230 192
rect 30 190 56 191
rect 95 190 165 191
rect 204 190 230 191
rect 30 189 57 190
rect 96 189 164 190
rect 203 189 230 190
rect 30 188 58 189
rect 97 188 163 189
rect 202 188 230 189
rect 30 187 59 188
rect 98 187 162 188
rect 201 187 230 188
rect 30 186 60 187
rect 99 186 161 187
rect 200 186 230 187
rect 30 185 61 186
rect 199 185 230 186
rect 30 184 62 185
rect 198 184 230 185
rect 30 183 63 184
rect 197 183 230 184
rect 30 182 64 183
rect 196 182 230 183
rect 30 181 65 182
rect 195 181 230 182
rect 30 180 66 181
rect 194 180 230 181
rect 30 179 67 180
rect 193 179 230 180
rect 30 178 68 179
rect 192 178 230 179
rect 30 177 69 178
rect 191 177 230 178
rect 30 176 70 177
rect 190 176 230 177
rect 30 175 71 176
rect 189 175 230 176
rect 30 174 72 175
rect 188 174 230 175
rect 30 173 73 174
rect 187 173 230 174
rect 30 172 74 173
rect 186 172 230 173
rect 30 171 75 172
rect 185 171 230 172
rect 30 170 76 171
rect 30 169 77 170
rect 30 168 78 169
rect 30 167 79 168
rect 30 105 80 167
rect 184 170 230 171
rect 183 169 230 170
rect 182 168 230 169
rect 181 167 230 168
rect 30 104 79 105
rect 30 103 78 104
rect 30 102 77 103
rect 30 101 76 102
rect 180 105 230 167
rect 181 104 230 105
rect 182 103 230 104
rect 183 102 230 103
rect 184 101 230 102
rect 30 100 75 101
rect 185 100 230 101
rect 30 99 74 100
rect 186 99 230 100
rect 30 98 73 99
rect 187 98 230 99
rect 30 97 72 98
rect 188 97 230 98
rect 30 96 71 97
rect 189 96 230 97
rect 30 95 70 96
rect 190 95 230 96
rect 30 94 69 95
rect 191 94 230 95
rect 30 93 68 94
rect 192 93 230 94
rect 30 92 67 93
rect 193 92 230 93
rect 30 91 66 92
rect 194 91 230 92
rect 30 90 65 91
rect 195 90 230 91
rect 30 89 64 90
rect 196 89 230 90
rect 30 88 63 89
rect 197 88 230 89
rect 30 87 62 88
rect 198 87 230 88
rect 30 86 61 87
rect 199 86 230 87
rect 30 85 60 86
rect 99 85 161 86
rect 200 85 230 86
rect 30 84 59 85
rect 98 84 162 85
rect 201 84 230 85
rect 30 83 58 84
rect 97 83 163 84
rect 202 83 230 84
rect 30 82 57 83
rect 96 82 164 83
rect 203 82 230 83
rect 30 81 56 82
rect 95 81 165 82
rect 204 81 230 82
rect 30 80 55 81
rect 94 80 166 81
rect 205 80 230 81
rect 30 79 54 80
rect 93 79 167 80
rect 206 79 230 80
rect 30 78 53 79
rect 92 78 168 79
rect 207 78 230 79
rect 30 77 52 78
rect 91 77 169 78
rect 208 77 230 78
rect 30 76 51 77
rect 90 76 170 77
rect 209 76 230 77
rect 30 75 50 76
rect 89 75 171 76
rect 210 75 230 76
rect 30 74 49 75
rect 88 74 172 75
rect 211 74 230 75
rect 30 73 48 74
rect 87 73 173 74
rect 212 73 230 74
rect 30 72 47 73
rect 86 72 174 73
rect 213 72 230 73
rect 30 71 46 72
rect 85 71 175 72
rect 214 71 230 72
rect 30 70 45 71
rect 84 70 176 71
rect 215 70 230 71
rect 30 69 44 70
rect 83 69 177 70
rect 216 69 230 70
rect 30 68 43 69
rect 82 68 178 69
rect 217 68 230 69
rect 30 67 42 68
rect 81 67 179 68
rect 218 67 230 68
rect 30 66 41 67
rect 80 66 180 67
rect 219 66 230 67
rect 30 65 40 66
rect 79 65 181 66
rect 220 65 230 66
rect 30 64 39 65
rect 78 64 182 65
rect 221 64 230 65
rect 30 63 38 64
rect 77 63 183 64
rect 222 63 230 64
rect 30 62 37 63
rect 76 62 184 63
rect 223 62 230 63
rect 30 61 36 62
rect 75 61 185 62
rect 224 61 230 62
rect 30 60 35 61
rect 74 60 186 61
rect 225 60 230 61
rect 30 59 34 60
rect 73 59 187 60
rect 226 59 230 60
rect 30 58 33 59
rect 72 58 188 59
rect 227 58 230 59
rect 30 57 32 58
rect 71 57 189 58
rect 228 57 230 58
rect 30 56 31 57
rect 70 56 190 57
rect 229 56 230 57
rect 69 55 191 56
rect 68 54 192 55
rect 67 53 193 54
rect 66 52 194 53
rect 65 51 195 52
rect 64 50 196 51
rect 63 49 197 50
rect 62 48 198 49
rect 61 47 199 48
rect 60 46 200 47
rect 59 45 201 46
rect 58 44 202 45
rect 57 43 203 44
rect 56 42 204 43
rect 55 41 205 42
rect 54 40 206 41
rect 53 39 207 40
rect 52 38 208 39
rect 51 37 209 38
rect 50 36 210 37
<< pdiffusionstop >>
rect 20 245 230 246
rect 20 244 229 245
rect 20 243 228 244
rect 20 242 227 243
rect 20 241 226 242
rect 20 240 225 241
rect 20 239 224 240
rect 20 238 223 239
rect 20 237 222 238
rect 20 236 221 237
rect 20 45 30 236
rect 239 235 240 236
rect 238 234 240 235
rect 237 233 240 234
rect 236 232 240 233
rect 235 231 240 232
rect 234 230 240 231
rect 233 229 240 230
rect 232 228 240 229
rect 231 227 240 228
rect 20 44 29 45
rect 20 43 28 44
rect 20 42 27 43
rect 20 41 26 42
rect 20 40 25 41
rect 20 39 24 40
rect 20 38 23 39
rect 20 37 22 38
rect 20 36 21 37
rect 230 36 240 227
rect 39 35 240 36
rect 38 34 240 35
rect 37 33 240 34
rect 36 32 240 33
rect 35 31 240 32
rect 34 30 240 31
rect 33 29 240 30
rect 32 28 240 29
rect 31 27 240 28
rect 30 26 240 27
<< glass >>
rect 95 146 120 171
rect 140 146 165 171
rect 95 101 120 126
rect 140 101 165 126
<< end >>
