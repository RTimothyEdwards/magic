magic
tech scmos
timestamp 616380303
<< polysilicon >>
rect 338 168 340 171
rect 344 165 346 167
rect 391 168 393 171
rect 385 165 387 167
rect 338 158 340 160
rect 357 156 359 160
rect 372 156 374 160
rect 391 158 393 160
rect 357 154 374 156
rect 357 153 359 154
rect 344 151 354 153
rect 344 146 346 151
rect 358 151 359 153
rect 344 140 346 143
rect 343 121 346 123
rect 349 121 351 123
rect 343 116 345 121
rect 365 114 367 154
rect 372 153 374 154
rect 372 151 373 153
rect 377 151 387 153
rect 385 146 387 151
rect 385 140 387 143
rect 380 121 382 123
rect 385 121 388 123
rect 386 116 388 121
rect 345 112 386 114
rect 340 103 342 111
rect 358 102 360 105
rect 371 102 373 105
rect 389 103 391 111
rect 351 96 353 98
rect 377 96 379 98
rect 358 92 360 93
rect 371 92 373 93
rect 358 86 360 87
rect 371 86 373 87
rect 351 83 353 85
rect 377 83 379 85
rect 339 69 341 78
rect 358 73 360 78
rect 371 73 373 78
rect 389 69 391 78
rect 342 59 344 64
rect 387 59 389 64
rect 342 57 346 59
rect 349 57 351 59
rect 380 57 382 59
rect 385 57 389 59
rect 344 37 346 39
rect 385 37 387 39
rect 344 29 346 34
rect 344 27 354 29
rect 338 20 340 22
rect 356 21 358 27
rect 372 27 373 29
rect 385 29 387 34
rect 377 27 387 29
rect 372 21 374 27
rect 391 21 393 23
rect 344 14 346 16
rect 338 11 340 13
rect 385 14 387 16
rect 391 11 393 13
<< ndiffusion >>
rect 335 165 338 168
rect 336 161 338 165
rect 335 160 338 161
rect 340 164 343 168
rect 346 167 361 170
rect 359 165 361 167
rect 371 167 385 170
rect 371 165 372 167
rect 346 164 357 165
rect 340 160 346 164
rect 350 160 357 164
rect 359 160 372 165
rect 374 164 385 165
rect 388 164 391 168
rect 374 160 381 164
rect 385 160 391 164
rect 393 160 396 168
rect 331 96 340 103
rect 342 99 349 103
rect 353 99 358 102
rect 342 98 351 99
rect 331 92 351 96
rect 355 93 358 99
rect 360 98 363 102
rect 368 98 371 102
rect 360 93 371 98
rect 373 99 377 102
rect 381 99 389 103
rect 373 93 376 99
rect 379 98 389 99
rect 391 99 397 103
rect 391 96 392 99
rect 379 95 392 96
rect 336 87 351 92
rect 331 85 351 87
rect 379 86 394 95
rect 331 78 339 85
rect 341 82 351 83
rect 355 82 358 86
rect 341 78 350 82
rect 354 78 358 82
rect 360 82 371 86
rect 360 78 363 82
rect 368 78 371 82
rect 373 82 376 86
rect 379 85 392 86
rect 379 82 389 83
rect 373 78 379 82
rect 383 78 389 82
rect 391 82 392 85
rect 391 78 397 82
rect 343 20 346 21
rect 335 13 338 20
rect 340 17 346 20
rect 350 17 356 21
rect 340 13 343 17
rect 346 16 356 17
rect 358 16 372 21
rect 374 17 381 21
rect 385 17 391 21
rect 374 16 385 17
rect 358 14 361 16
rect 346 12 361 14
rect 371 14 372 16
rect 371 12 385 14
rect 388 13 391 17
rect 393 13 396 21
rect 346 11 385 12
<< pdiffusion >>
rect 339 143 344 146
rect 346 143 347 146
rect 339 139 343 143
rect 339 135 346 139
rect 339 128 347 135
rect 339 124 346 128
rect 346 123 349 124
rect 346 120 349 121
rect 346 117 354 120
rect 384 143 385 146
rect 387 143 392 146
rect 388 139 392 143
rect 385 135 392 139
rect 384 128 392 135
rect 385 124 392 128
rect 382 123 385 124
rect 382 120 385 121
rect 377 117 385 120
rect 346 60 354 63
rect 346 59 349 60
rect 377 60 385 63
rect 382 59 385 60
rect 346 56 349 57
rect 382 56 385 57
rect 339 52 346 56
rect 385 52 392 56
rect 339 45 347 52
rect 384 45 392 52
rect 339 41 346 45
rect 385 41 392 45
rect 339 37 343 41
rect 388 37 392 41
rect 339 34 344 37
rect 346 34 347 37
rect 384 34 385 37
rect 387 34 392 37
<< metal1 >>
rect 339 176 342 178
rect 341 171 342 176
rect 331 159 336 161
rect 339 152 342 171
rect 334 149 342 152
rect 334 106 337 149
rect 347 147 350 160
rect 354 160 357 178
rect 366 171 367 176
rect 366 170 371 171
rect 374 160 377 178
rect 389 176 392 178
rect 389 171 390 176
rect 354 156 364 160
rect 340 143 347 146
rect 340 116 343 143
rect 346 134 350 135
rect 346 129 348 134
rect 346 128 350 129
rect 355 121 358 148
rect 350 117 354 120
rect 334 103 346 106
rect 350 103 353 117
rect 361 114 364 156
rect 343 75 346 103
rect 357 111 364 114
rect 367 156 377 160
rect 367 114 370 156
rect 373 121 376 148
rect 381 147 384 160
rect 389 152 392 171
rect 389 149 397 152
rect 384 143 391 146
rect 381 134 385 135
rect 383 129 385 134
rect 381 128 385 129
rect 367 111 374 114
rect 357 92 360 111
rect 363 102 368 104
rect 371 92 374 111
rect 377 103 380 120
rect 388 116 391 143
rect 394 106 397 149
rect 386 103 397 106
rect 357 87 358 92
rect 373 87 374 92
rect 333 72 346 75
rect 333 31 336 72
rect 339 37 343 64
rect 351 60 354 78
rect 357 69 360 87
rect 363 76 368 78
rect 371 69 374 87
rect 357 66 364 69
rect 346 51 350 52
rect 346 46 348 51
rect 346 45 350 46
rect 339 34 347 37
rect 333 28 342 31
rect 331 19 335 21
rect 339 11 342 28
rect 347 21 350 33
rect 355 32 358 59
rect 361 24 364 66
rect 354 21 364 24
rect 367 66 374 69
rect 367 24 370 66
rect 379 63 382 78
rect 386 75 389 103
rect 392 92 399 95
rect 392 87 395 92
rect 392 86 399 87
rect 386 72 398 75
rect 377 60 382 63
rect 373 32 376 59
rect 381 51 385 52
rect 383 46 385 51
rect 381 45 385 46
rect 388 37 392 64
rect 384 34 392 37
rect 367 21 377 24
rect 341 6 342 11
rect 339 4 342 6
rect 354 4 357 21
rect 361 11 371 12
rect 365 10 371 11
rect 365 6 366 10
rect 374 4 377 21
rect 381 21 384 33
rect 395 31 398 72
rect 389 28 398 31
rect 389 11 392 28
rect 389 6 390 11
rect 389 4 392 6
<< metal2 >>
rect 331 171 367 176
rect 371 171 402 176
rect 331 154 336 155
rect 331 150 402 154
rect 331 129 348 134
rect 352 129 379 134
rect 383 129 402 134
rect 331 119 402 123
rect 331 110 402 114
rect 363 108 368 110
rect 331 87 395 92
rect 399 87 402 92
rect 363 70 368 72
rect 331 66 402 70
rect 331 57 402 61
rect 331 46 348 51
rect 352 46 379 51
rect 383 46 402 51
rect 331 26 402 30
rect 331 25 336 26
rect 331 10 402 11
rect 331 6 366 10
rect 371 6 402 10
<< polycontact >>
rect 336 171 341 176
rect 390 171 395 176
rect 354 148 358 153
rect 340 111 345 116
rect 373 148 377 153
rect 386 111 391 116
rect 358 87 363 92
rect 368 87 373 92
rect 339 64 344 69
rect 387 64 392 69
rect 354 27 358 32
rect 373 27 377 32
rect 336 6 341 11
rect 390 6 395 11
<< ndcontact >>
rect 331 161 336 165
rect 361 165 371 170
rect 346 160 350 164
rect 381 160 385 164
rect 349 99 353 103
rect 363 98 368 102
rect 377 99 381 103
rect 392 95 402 99
rect 350 78 354 82
rect 363 78 368 82
rect 379 78 383 82
rect 392 82 402 86
rect 331 15 335 19
rect 346 17 350 21
rect 381 17 385 21
rect 361 12 371 16
<< pdcontact >>
rect 347 143 351 147
rect 346 124 350 128
rect 354 117 358 121
rect 380 143 384 147
rect 381 124 385 128
rect 373 117 377 121
rect 354 59 358 63
rect 373 59 377 63
rect 346 52 350 56
rect 381 52 385 56
rect 347 33 351 37
rect 380 33 384 37
<< m2contact >>
rect 331 155 336 159
rect 367 171 371 176
rect 348 129 352 134
rect 379 129 383 134
rect 363 104 368 108
rect 363 72 368 76
rect 348 46 352 51
rect 331 21 335 25
rect 395 87 399 92
rect 379 46 383 51
rect 366 6 371 10
<< ntransistor >>
rect 338 160 340 168
rect 346 165 359 167
rect 372 165 385 167
rect 357 160 359 165
rect 372 160 374 165
rect 391 160 393 168
rect 340 98 342 103
rect 340 96 351 98
rect 358 93 360 102
rect 371 93 373 102
rect 389 98 391 103
rect 379 96 391 98
rect 339 83 351 85
rect 339 78 341 83
rect 358 78 360 86
rect 371 78 373 86
rect 379 83 391 85
rect 389 78 391 83
rect 338 13 340 20
rect 356 16 358 21
rect 372 16 374 21
rect 346 14 358 16
rect 372 14 385 16
rect 391 13 393 21
<< ptransistor >>
rect 344 143 346 146
rect 346 121 349 123
rect 385 143 387 146
rect 382 121 385 123
rect 346 57 349 59
rect 382 57 385 59
rect 344 34 346 37
rect 385 34 387 37
<< psubstratepcontact >>
rect 361 170 366 176
rect 331 87 336 92
rect 361 6 365 11
<< nsubstratencontact >>
rect 346 135 350 139
rect 381 135 385 139
rect 346 41 350 45
rect 381 41 385 45
<< labels >>
rlabel metal2 402 89 402 89 7 GND!
rlabel metal1 391 178 391 178 5 accA1#
rlabel metal1 355 178 355 178 5 accB0#
rlabel metal1 376 178 376 178 5 accB1#
rlabel metal1 340 178 340 178 5 accA0#
rlabel space 359 125 378 143 5 Plow here
rlabel metal2 402 112 402 112 7 busB1#
rlabel metal2 402 68 402 68 7 busB0#
rlabel metal2 402 49 402 49 7 Vdd!
rlabel metal2 402 28 402 28 7 busA0#
rlabel metal1 391 4 391 4 1 accA1#
rlabel metal1 340 4 340 4 1 accA0#
rlabel metal2 402 9 402 9 8 GND!
rlabel metal1 355 4 355 4 1 accB0#
rlabel metal1 376 4 376 4 1 accB1#
<< end >>
