magic
tech scmos
timestamp 955571370
<< error_p >>
rect 22 21 26 25
rect 22 16 26 18
rect 22 12 26 15
rect 22 10 26 11
rect 21 6 22 10
rect 26 6 27 10
rect 22 5 26 6
rect 21 1 22 5
rect 26 1 27 5
rect 22 0 26 1
<< polysilicon >>
rect 1 30 6 32
rect 9 30 13 32
rect 22 26 26 30
rect 1 6 6 8
rect 9 6 12 8
<< ndiffusion >>
rect 22 16 26 20
rect 6 8 9 10
rect 6 4 9 6
<< pdiffusion >>
rect 6 32 9 33
rect 6 29 9 30
rect 22 21 26 25
<< metal1 >>
rect 1 34 6 37
rect 10 34 15 37
rect 22 31 26 35
rect 6 22 10 25
rect 6 18 15 22
rect 6 14 10 18
rect 1 0 6 3
rect 10 0 15 3
<< ntransistor >>
rect 6 6 9 8
rect 22 1 26 5
<< ptransistor >>
rect 6 30 9 32
rect 22 6 26 10
<< ndcontact >>
rect 6 10 10 14
rect 22 11 26 15
rect 6 0 10 4
<< pdcontact >>
rect 6 33 10 37
rect 6 25 10 29
<< labels >>
rlabel metal1 22 31 26 35 3 Metal
rlabel polysilicon 22 26 26 30 3 Polysilicon
rlabel pdiffusion 22 21 26 25 3 P-Diffusion
rlabel ndiffusion 22 16 26 20 3 N-Diffusion
rlabel ndcontact 22 11 26 15 3 Contact
rlabel ptransistor 22 6 26 10 3 P-Fet
rlabel ntransistor 22 1 26 5 3 N-Fet
<< end >>
