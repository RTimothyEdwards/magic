magic
tech scmos
timestamp 760840608
<< polysilicon >>
rect 383 99 398 102
rect 383 98 385 99
rect 356 95 385 98
rect 389 95 391 99
rect 395 95 398 99
rect 356 94 398 95
rect 356 92 360 94
rect 356 88 390 92
rect 386 85 390 88
rect 356 81 390 85
rect 356 78 360 81
rect 356 74 390 78
rect 386 72 390 74
rect 356 68 390 72
rect 356 66 360 68
rect 356 62 390 66
rect 386 59 390 62
rect 356 55 390 59
rect 356 52 360 55
rect 356 51 398 52
rect 356 48 385 51
rect 383 47 385 48
rect 389 47 391 51
rect 395 47 398 51
rect 383 45 398 47
<< metal1 >>
rect 446 152 453 153
rect 445 151 453 152
rect 444 150 453 151
rect 443 149 453 150
rect 442 148 453 149
rect 441 147 453 148
rect 440 146 452 147
rect 439 145 451 146
rect 438 144 450 145
rect 437 143 449 144
rect 436 142 448 143
rect 435 141 447 142
rect 434 140 446 141
rect 433 139 445 140
rect 432 138 444 139
rect 431 137 443 138
rect 430 136 442 137
rect 429 135 441 136
rect 428 134 440 135
rect 427 133 439 134
rect 426 132 438 133
rect 425 131 437 132
rect 424 130 436 131
rect 423 129 435 130
rect 422 128 434 129
rect 421 127 433 128
rect 420 126 432 127
rect 419 125 431 126
rect 418 124 430 125
rect 417 123 429 124
rect 416 122 428 123
rect 415 121 427 122
rect 414 120 426 121
rect 413 119 425 120
rect 412 118 424 119
rect 411 117 423 118
rect 410 116 422 117
rect 409 115 421 116
rect 408 114 420 115
rect 407 113 419 114
rect 406 112 418 113
rect 405 111 417 112
rect 404 110 416 111
rect 403 109 415 110
rect 402 108 414 109
rect 401 107 413 108
rect 400 106 412 107
rect 399 105 411 106
rect 398 104 410 105
rect 397 103 409 104
rect 396 102 408 103
rect 383 101 407 102
rect 383 100 406 101
rect 383 99 405 100
rect 383 95 385 99
rect 389 95 391 99
rect 395 98 404 99
rect 395 97 403 98
rect 395 96 402 97
rect 395 95 401 96
rect 383 94 400 95
rect 383 93 399 94
rect 383 52 402 53
rect 383 51 403 52
rect 383 47 385 51
rect 389 47 391 51
rect 395 50 404 51
rect 395 49 405 50
rect 395 48 406 49
rect 395 47 407 48
rect 383 46 408 47
rect 383 45 409 46
rect 396 44 410 45
rect 397 43 411 44
rect 398 42 412 43
rect 399 41 413 42
rect 400 40 414 41
rect 401 39 415 40
rect 402 38 416 39
rect 403 37 417 38
rect 404 36 418 37
rect 405 35 419 36
rect 406 34 420 35
rect 407 33 421 34
rect 408 32 422 33
rect 409 31 423 32
rect 410 30 424 31
rect 411 29 425 30
rect 412 28 426 29
rect 413 27 427 28
rect 414 26 428 27
rect 415 25 429 26
rect 416 24 430 25
rect 417 23 431 24
rect 418 22 432 23
rect 419 21 433 22
rect 420 20 434 21
rect 421 19 435 20
rect 422 18 436 19
rect 423 17 437 18
rect 424 16 438 17
rect 425 15 439 16
rect 426 14 440 15
rect 427 13 441 14
rect 428 12 442 13
rect 429 11 443 12
rect 430 10 444 11
rect 431 9 445 10
rect 432 8 446 9
rect 433 7 447 8
rect 434 6 448 7
rect 435 5 449 6
rect 436 4 450 5
rect 437 3 451 4
rect 438 2 452 3
rect 439 1 453 2
rect 440 0 453 1
rect 441 -1 453 0
rect 442 -2 453 -1
rect 443 -3 453 -2
rect 444 -4 453 -3
rect 445 -5 453 -4
rect 446 -6 453 -5
rect 447 -7 453 -6
<< polycontact >>
rect 385 95 389 99
rect 391 95 395 99
rect 385 47 389 51
rect 391 47 395 51
<< substrateopen >>
rect 309 152 438 153
rect 310 151 437 152
rect 311 150 436 151
rect 312 149 435 150
rect 313 148 434 149
rect 314 147 433 148
rect 315 146 432 147
rect 316 145 431 146
rect 317 144 430 145
rect 318 143 429 144
rect 319 142 428 143
rect 320 141 427 142
rect 321 140 426 141
rect 322 139 425 140
rect 293 138 294 139
rect 323 138 424 139
rect 452 138 453 139
rect 293 137 295 138
rect 324 137 423 138
rect 451 137 453 138
rect 293 136 296 137
rect 325 136 422 137
rect 450 136 453 137
rect 293 135 297 136
rect 326 135 421 136
rect 449 135 453 136
rect 293 134 298 135
rect 327 134 420 135
rect 448 134 453 135
rect 293 133 299 134
rect 328 133 419 134
rect 447 133 453 134
rect 293 132 300 133
rect 329 132 418 133
rect 446 132 453 133
rect 293 131 301 132
rect 330 131 417 132
rect 445 131 453 132
rect 293 130 302 131
rect 331 130 416 131
rect 444 130 453 131
rect 293 129 303 130
rect 332 129 415 130
rect 443 129 453 130
rect 293 128 304 129
rect 333 128 414 129
rect 442 128 453 129
rect 293 127 305 128
rect 334 127 413 128
rect 441 127 453 128
rect 293 126 306 127
rect 335 126 412 127
rect 440 126 453 127
rect 293 125 307 126
rect 336 125 411 126
rect 439 125 453 126
rect 293 124 308 125
rect 337 124 410 125
rect 438 124 453 125
rect 293 123 309 124
rect 338 123 409 124
rect 437 123 453 124
rect 293 122 310 123
rect 339 122 408 123
rect 436 122 453 123
rect 293 121 311 122
rect 340 121 407 122
rect 435 121 453 122
rect 293 120 312 121
rect 341 120 406 121
rect 434 120 453 121
rect 293 119 313 120
rect 342 119 405 120
rect 433 119 453 120
rect 293 118 314 119
rect 343 118 404 119
rect 432 118 453 119
rect 293 117 315 118
rect 344 117 403 118
rect 431 117 453 118
rect 293 116 316 117
rect 345 116 402 117
rect 430 116 453 117
rect 293 115 317 116
rect 346 115 401 116
rect 429 115 453 116
rect 293 114 318 115
rect 347 114 400 115
rect 428 114 453 115
rect 293 113 319 114
rect 348 113 399 114
rect 427 113 453 114
rect 293 112 320 113
rect 349 112 398 113
rect 426 112 453 113
rect 293 111 321 112
rect 350 111 397 112
rect 425 111 453 112
rect 293 110 322 111
rect 351 110 396 111
rect 424 110 453 111
rect 293 109 323 110
rect 352 109 395 110
rect 423 109 453 110
rect 293 108 324 109
rect 353 108 394 109
rect 422 108 453 109
rect 293 107 325 108
rect 354 107 393 108
rect 421 107 453 108
rect 293 106 326 107
rect 355 106 392 107
rect 420 106 453 107
rect 293 105 327 106
rect 356 105 391 106
rect 419 105 453 106
rect 293 104 328 105
rect 418 104 453 105
rect 293 103 329 104
rect 417 103 453 104
rect 293 102 330 103
rect 416 102 453 103
rect 293 101 331 102
rect 415 101 453 102
rect 293 100 332 101
rect 414 100 453 101
rect 293 99 333 100
rect 413 99 453 100
rect 293 98 334 99
rect 412 98 453 99
rect 293 97 335 98
rect 411 97 453 98
rect 293 96 336 97
rect 410 96 453 97
rect 293 95 337 96
rect 409 95 453 96
rect 293 94 338 95
rect 408 94 453 95
rect 293 93 339 94
rect 407 93 453 94
rect 293 92 340 93
rect 406 92 453 93
rect 293 57 341 92
rect 405 57 453 92
rect 293 56 340 57
rect 406 56 453 57
rect 293 55 339 56
rect 407 55 453 56
rect 293 54 338 55
rect 408 54 453 55
rect 293 53 337 54
rect 409 53 453 54
rect 293 52 336 53
rect 410 52 453 53
rect 293 51 335 52
rect 411 51 453 52
rect 293 50 334 51
rect 412 50 453 51
rect 293 49 333 50
rect 413 49 453 50
rect 293 48 332 49
rect 414 48 453 49
rect 293 47 331 48
rect 415 47 453 48
rect 293 46 330 47
rect 416 46 453 47
rect 293 45 329 46
rect 417 45 453 46
rect 293 44 328 45
rect 418 44 453 45
rect 293 43 327 44
rect 419 43 453 44
rect 293 42 326 43
rect 420 42 453 43
rect 293 41 325 42
rect 421 41 453 42
rect 293 40 324 41
rect 356 40 391 41
rect 422 40 453 41
rect 293 39 323 40
rect 355 39 392 40
rect 423 39 453 40
rect 293 38 322 39
rect 354 38 393 39
rect 424 38 453 39
rect 293 37 321 38
rect 353 37 394 38
rect 425 37 453 38
rect 293 36 320 37
rect 352 36 395 37
rect 426 36 453 37
rect 293 35 319 36
rect 351 35 396 36
rect 427 35 453 36
rect 293 34 318 35
rect 350 34 397 35
rect 428 34 453 35
rect 293 33 317 34
rect 349 33 398 34
rect 429 33 453 34
rect 293 32 316 33
rect 348 32 399 33
rect 430 32 453 33
rect 293 31 315 32
rect 347 31 400 32
rect 431 31 453 32
rect 293 30 314 31
rect 346 30 401 31
rect 432 30 453 31
rect 293 29 313 30
rect 345 29 402 30
rect 433 29 453 30
rect 293 28 312 29
rect 344 28 403 29
rect 434 28 453 29
rect 293 27 311 28
rect 343 27 404 28
rect 435 27 453 28
rect 293 26 310 27
rect 342 26 405 27
rect 436 26 453 27
rect 293 25 309 26
rect 341 25 406 26
rect 437 25 453 26
rect 293 24 308 25
rect 340 24 407 25
rect 438 24 453 25
rect 293 23 307 24
rect 339 23 408 24
rect 439 23 453 24
rect 293 22 306 23
rect 338 22 409 23
rect 440 22 453 23
rect 293 21 305 22
rect 337 21 410 22
rect 441 21 453 22
rect 293 20 304 21
rect 336 20 411 21
rect 442 20 453 21
rect 293 19 303 20
rect 335 19 412 20
rect 443 19 453 20
rect 293 18 302 19
rect 334 18 413 19
rect 444 18 453 19
rect 293 17 301 18
rect 333 17 414 18
rect 445 17 453 18
rect 293 16 300 17
rect 332 16 415 17
rect 446 16 453 17
rect 293 15 299 16
rect 331 15 416 16
rect 447 15 453 16
rect 293 14 298 15
rect 330 14 417 15
rect 448 14 453 15
rect 293 13 297 14
rect 329 13 418 14
rect 449 13 453 14
rect 293 12 296 13
rect 328 12 419 13
rect 450 12 453 13
rect 293 11 295 12
rect 327 11 420 12
rect 451 11 453 12
rect 293 10 294 11
rect 326 10 421 11
rect 452 10 453 11
rect 325 9 422 10
rect 324 8 423 9
rect 323 7 424 8
rect 322 6 425 7
rect 321 5 426 6
rect 320 4 427 5
rect 319 3 428 4
rect 318 2 429 3
rect 317 1 430 2
rect 316 0 431 1
rect 315 -1 432 0
rect 314 -2 433 -1
rect 313 -3 434 -2
rect 312 -4 435 -3
rect 311 -5 436 -4
rect 310 -6 437 -5
rect 309 -7 438 -6
<< pdiffusionstop >>
rect 288 153 458 158
rect 288 -7 293 153
rect 453 -7 458 153
rect 288 -12 458 -7
<< end >>
