magic
tech scmos
timestamp 736070890
<< nwell >>
rect -2 -2 20 8
<< ndiffusion >>
rect 0 13 4 16
rect 7 13 11 16
<< pdiffusion >>
rect 0 0 4 3
rect 7 0 11 3
<< psubstratepdiff >>
rect 15 11 18 16
<< nsubstratendiff >>
rect 15 0 18 5
<< labels >>
rlabel nwell -1 8 20 8 1 P-Region
rlabel nwell -1 8 20 8 5 N-Region
rlabel space -1 13 -1 16 3 2.1
rlabel space 4 12 7 12 1 2.2
rlabel space 17 8 17 11 3 2.4
rlabel space 12 8 12 13 3 2.3
rlabel nwell 6 3 6 8 3 2.3
<< end >>
