magic
tech scmos
timestamp 736115372
<< capwell >>
rect -3 -3 129 122
<< polysilicon >>
rect -1 103 0 107
rect -1 80 0 84
rect -1 57 0 61
rect -1 34 0 38
rect -1 11 0 15
<< wellcapacitor >>
rect 3 107 23 115
rect 26 107 46 115
rect 49 107 69 115
rect 72 107 92 115
rect 95 107 115 115
rect 3 103 115 107
rect 3 95 23 103
rect 26 95 46 103
rect 49 95 69 103
rect 72 95 92 103
rect 95 95 115 103
rect 11 92 15 95
rect 34 92 38 95
rect 57 92 61 95
rect 80 92 84 95
rect 103 92 107 95
rect 3 84 23 92
rect 26 84 46 92
rect 49 84 69 92
rect 72 84 92 92
rect 95 84 115 92
rect 3 80 115 84
rect 3 72 23 80
rect 26 72 46 80
rect 49 72 69 80
rect 72 72 92 80
rect 95 72 115 80
rect 11 69 15 72
rect 34 69 38 72
rect 57 69 61 72
rect 80 69 84 72
rect 103 69 107 72
rect 3 61 23 69
rect 26 61 46 69
rect 49 61 69 69
rect 72 61 92 69
rect 95 61 115 69
rect 3 57 115 61
rect 3 49 23 57
rect 26 49 46 57
rect 49 49 69 57
rect 72 49 92 57
rect 95 49 115 57
rect 11 46 15 49
rect 34 46 38 49
rect 57 46 61 49
rect 80 46 84 49
rect 103 46 107 49
rect 3 38 23 46
rect 26 38 46 46
rect 49 38 69 46
rect 72 38 92 46
rect 95 38 115 46
rect 3 34 115 38
rect 3 26 23 34
rect 26 26 46 34
rect 49 26 69 34
rect 72 26 92 34
rect 95 26 115 34
rect 11 23 15 26
rect 34 23 38 26
rect 57 23 61 26
rect 80 23 84 26
rect 103 23 107 26
rect 3 15 23 23
rect 26 15 46 23
rect 49 15 69 23
rect 72 15 92 23
rect 95 15 115 23
rect 3 11 115 15
rect 3 3 23 11
rect 26 3 46 11
rect 49 3 69 11
rect 72 3 92 11
rect 95 3 115 11
<< ndiffusion >>
rect 0 115 119 119
rect 0 107 3 115
rect 23 107 26 115
rect 46 107 49 115
rect 69 107 72 115
rect 92 107 95 115
rect 0 95 3 103
rect 23 95 26 103
rect 46 95 49 103
rect 69 95 72 103
rect 92 95 95 103
rect 115 95 119 115
rect 0 92 11 95
rect 15 92 34 95
rect 38 92 57 95
rect 61 92 80 95
rect 84 92 103 95
rect 107 92 119 95
rect 0 84 3 92
rect 23 84 26 92
rect 46 84 49 92
rect 69 84 72 92
rect 92 84 95 92
rect 0 72 3 80
rect 23 72 26 80
rect 46 72 49 80
rect 69 72 72 80
rect 92 72 95 80
rect 115 72 119 92
rect 0 69 11 72
rect 15 69 34 72
rect 38 69 57 72
rect 61 69 80 72
rect 84 69 103 72
rect 107 69 119 72
rect 0 61 3 69
rect 23 61 26 69
rect 46 61 49 69
rect 69 61 72 69
rect 92 61 95 69
rect 0 49 3 57
rect 23 49 26 57
rect 46 49 49 57
rect 69 49 72 57
rect 92 49 95 57
rect 115 49 119 69
rect 0 46 11 49
rect 15 46 34 49
rect 38 46 57 49
rect 61 46 80 49
rect 84 46 103 49
rect 107 46 119 49
rect 0 38 3 46
rect 23 38 26 46
rect 46 38 49 46
rect 69 38 72 46
rect 92 38 95 46
rect 0 26 3 34
rect 23 26 26 34
rect 46 26 49 34
rect 69 26 72 34
rect 92 26 95 34
rect 115 26 119 46
rect 0 23 11 26
rect 15 23 34 26
rect 38 23 57 26
rect 61 23 80 26
rect 84 23 103 26
rect 107 23 119 26
rect 0 15 3 23
rect 23 15 26 23
rect 46 15 49 23
rect 69 15 72 23
rect 92 15 95 23
rect 0 3 3 11
rect 23 3 26 11
rect 46 3 49 11
rect 69 3 72 11
rect 92 3 95 11
rect 115 3 119 23
rect 0 0 119 3
<< ntransistor >>
rect 0 103 3 107
rect 0 80 3 84
rect 0 57 3 61
rect 0 34 3 38
rect 0 11 3 15
<< polycontact >>
rect -5 3 -1 115
<< ndcontact >>
rect 119 0 123 119
<< end >>
