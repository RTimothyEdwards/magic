magic
tech scmos
timestamp 801256319
<< nwell >>
rect 0 -1 20 13
<< metal1 >>
rect -1 4 5 8
rect 17 4 21 8
<< pdcontact >>
rect 5 4 9 8
<< psubstratepcontact >>
rect -7 16 27 20
rect -7 -8 27 -4
<< nsubstratencontact >>
rect 13 4 17 8
<< psubstratepdiff >>
rect -7 -4 -3 16
rect 23 -4 27 16
<< labels >>
rlabel metal1 21 6 21 6 3 base
rlabel metal1 -1 6 -1 6 7 emitter
rlabel psubstratepcontact 10 18 10 18 1 collector
rlabel psubstratepcontact 10 -6 10 -6 5 collector
<< end >>
