magic
tech scmos
timestamp 500615676
<< polysilicon >>
rect 4 2 6 10
rect 4 -5 6 -1
rect 4 -15 6 -8
<< ndiffusion >>
rect -5 -1 4 2
rect 6 -1 8 2
rect -5 -8 4 -5
rect 6 -8 8 -5
<< metal1 >>
rect -7 11 2 14
rect 7 11 30 14
<< polycontact >>
rect 2 10 7 14
<< ntransistor >>
rect 4 -1 6 2
rect 4 -8 6 -5
<< labels >>
rlabel metal1 24 12 24 12 1 Local node name
rlabel ndiffusion -3 -6 -3 -6 1 Global name!
rlabel ndiffusion -3 1 -3 1 1 Node Attribute@
rlabel ntransistor 6 1 6 1 3 Source/Drain Attribute$
rlabel ntransistor 5 -6 5 -6 3 Gate Attribute^
rlabel metal1 -7 11 -7 14 7 Label for routing
<< end >>
