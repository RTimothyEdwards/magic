magic
tech scmos
timestamp 617322824
<< polysilicon >>
rect -13 8 -9 10
rect -6 8 10 10
rect -13 1 -9 5
rect -6 1 -3 5
<< ndiffusion >>
rect -9 10 -6 13
rect -9 5 -6 8
rect -9 -1 -6 1
rect -9 -9 -6 -5
<< metal1 >>
rect 1 1 10 4
rect -6 -5 10 -2
<< polycontact >>
rect -3 1 1 5
<< ndcontact >>
rect -10 -5 -6 -1
<< ntransistor >>
rect -9 8 -6 10
rect -9 1 -6 5
<< end >>
