magic
tech scmos
timestamp 539497029
<< metal1 >>
rect -6 24 4 28
rect -40 -3 -36 4
rect -6 -22 -2 24
rect 1 -3 5 4
rect 5 -7 24 -3
rect -6 -26 4 -22
<< metal2 >>
rect -36 -7 1 -4
<< m2contact >>
rect -40 -7 -36 -3
rect 1 -7 5 -3
<< labels >>
rlabel metal1 24 -5 24 -5 3 ReceiverC
rlabel metal1 3 4 3 4 1 Driver2
rlabel metal1 -38 4 -38 4 1 ReceiverB
rlabel metal1 4 -24 4 -24 3 Driver1
rlabel metal1 4 27 4 27 3 ReceiverA
<< end >>
