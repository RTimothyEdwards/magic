magic
tech scmos
timestamp 796597909
<< nwell >>
rect -28 -20 30 38
<< metal1 >>
rect -38 41 -35 45
rect 32 41 33 45
rect -38 30 -23 34
rect 21 33 26 34
rect 21 30 22 33
rect -8 18 -6 22
rect 8 21 14 22
rect 8 18 10 21
rect -38 7 -1 11
rect -38 -4 -12 0
rect -8 -4 -6 0
rect 8 -3 10 0
rect 8 -4 14 -3
rect 21 -15 22 -12
rect 21 -16 26 -15
rect -38 -27 -35 -23
rect 32 -27 33 -23
<< collector >>
rect -25 34 27 35
rect -25 30 -23 34
rect 21 33 27 34
rect 21 30 22 33
rect -25 29 22 30
rect -25 -11 -19 29
rect 21 -11 22 29
rect -25 -12 22 -11
rect -25 -16 -23 -12
rect 21 -15 22 -12
rect 26 -15 27 33
rect 21 -16 27 -15
rect -25 -17 27 -16
<< pbase >>
rect -15 22 17 25
rect -15 14 -12 22
rect -8 18 -6 22
rect 8 21 17 22
rect 8 18 10 21
rect -8 14 10 18
rect -15 11 10 14
rect -15 7 -1 11
rect 3 7 10 11
rect -15 4 10 7
rect -15 -4 -12 4
rect -8 0 10 4
rect -8 -4 -6 0
rect 8 -3 10 0
rect 14 -3 17 21
rect 8 -4 17 -3
rect -15 -7 17 -4
<< collectorcontact >>
rect -23 30 21 34
rect -23 -16 21 -12
rect 22 -15 26 33
<< emittercontact >>
rect -1 7 3 11
<< pbasecontact >>
rect -12 14 -8 22
rect -6 18 8 22
rect -12 -4 -8 4
rect -6 -4 8 0
rect 10 -3 14 21
<< psubstratepcontact >>
rect -35 41 32 45
rect -35 -27 32 -23
rect 33 -27 37 45
<< psubstratepdiff >>
rect 32 41 33 45
rect -35 -23 -31 41
rect 32 -27 33 -23
<< labels >>
rlabel metal1 -37 9 -37 9 4 EMITTER
rlabel metal1 -37 -2 -37 -2 2 BASE
rlabel metal1 -37 -25 -37 -25 2 GUARDRING
rlabel metal1 -37 43 -37 43 4 GND
rlabel metal1 -37 32 -37 32 4 COLLECTOR
<< end >>
