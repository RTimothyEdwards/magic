magic
tech scmos
timestamp 715648344
<< polysilicon >>
rect 11 0 13 6
<< ndiffusion >>
rect 2 4 5 11
<< metal1 >>
rect 0 7 10 10
rect 5 0 15 3
<< polycontact >>
rect 10 6 14 10
<< ndcontact >>
rect 1 0 5 4
<< labels >>
rlabel space 0 3 0 4 7 7.4
rlabel space 17 0 17 3 3 7.1
rlabel space 15 6 15 7 3 7.3
rlabel space 18 3 18 6 3 7.2
<< end >>
