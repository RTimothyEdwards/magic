magic
tech scmos
timestamp 617565736
<< polysilicon >>
rect -95 26 -92 28
rect -72 26 -70 28
rect -3 26 0 28
rect 4 26 6 28
rect -95 2 -93 26
rect -3 17 -1 26
rect -72 15 -1 17
rect -3 2 -1 15
rect -95 0 -92 2
rect -72 0 -70 2
rect -3 0 0 2
rect 4 0 8 2
rect 6 -16 8 0
rect -95 -18 -92 -16
rect -72 -18 -70 -16
rect -2 -18 0 -16
rect 4 -18 18 -16
rect -95 -42 -93 -18
rect -3 -22 0 -20
rect 4 -22 6 -20
rect -3 -31 -1 -22
rect -72 -33 -1 -31
rect -3 -42 -1 -33
rect 16 -42 18 -18
rect -95 -44 -92 -42
rect -72 -44 -70 -42
rect -3 -44 0 -42
rect 4 -44 6 -42
rect 8 -44 10 -42
rect 14 -44 18 -42
<< ndiffusion >>
rect -92 2 -72 3
rect 0 2 4 3
rect -92 -1 -72 0
rect 0 -1 4 0
rect -92 -16 -72 -15
rect 0 -16 4 -15
rect -92 -19 -72 -18
rect 0 -20 4 -18
rect 0 -23 4 -22
<< pdiffusion >>
rect -92 28 -72 29
rect 0 28 4 29
rect -92 25 -72 26
rect 0 25 4 26
rect -92 -42 -72 -41
rect 0 -42 4 -41
rect 10 -42 14 -41
rect -92 -45 -72 -44
rect 0 -45 4 -44
rect 10 -45 14 -44
<< metal1 >>
rect -88 34 -87 38
rect -92 33 -87 34
rect -1 34 0 38
rect -5 33 0 34
rect -76 18 -72 21
rect -102 14 -99 18
rect -76 7 -72 14
rect 0 7 4 21
rect -92 -6 -87 -5
rect -88 -10 -87 -6
rect -92 -11 -87 -10
rect -5 -6 0 -5
rect -1 -10 0 -6
rect -5 -11 0 -10
rect -76 -30 -72 -23
rect -103 -34 -99 -30
rect -76 -37 -72 -34
rect 0 -37 4 -27
rect 4 -41 10 -37
rect 4 -49 10 -45
rect -92 -50 -87 -49
rect -88 -54 -87 -50
rect -5 -50 0 -49
rect -1 -54 0 -50
<< metal2 >>
rect -104 34 -92 38
rect -88 34 -5 38
rect -1 34 24 38
rect 20 -6 24 34
rect -110 -10 -92 -6
rect -88 -10 -5 -6
rect -1 -10 13 -6
rect 20 -10 28 -6
rect 20 -50 24 -10
rect -104 -54 -92 -50
rect -88 -54 -5 -50
rect -1 -54 24 -50
<< nwell >>
rect -101 16 -70 39
rect -14 16 17 39
rect -101 -55 -70 -32
rect -14 -55 17 -32
<< polycontact >>
rect -99 14 -95 18
rect -76 14 -72 18
rect -99 -34 -95 -30
rect -76 -34 -72 -30
<< ndcontact >>
rect -92 3 -72 7
rect 0 3 4 7
rect -92 -5 -72 -1
rect 0 -5 4 -1
rect -92 -15 -72 -11
rect 0 -15 4 -11
rect -92 -23 -72 -19
rect 0 -27 4 -23
<< pdcontact >>
rect -92 29 -72 33
rect 0 29 4 33
rect -92 21 -72 25
rect 0 21 4 25
rect -92 -41 -72 -37
rect 0 -41 4 -37
rect 10 -41 14 -37
rect -92 -49 -72 -45
rect 0 -49 4 -45
rect 10 -49 14 -45
<< m2contact >>
rect -92 34 -88 38
rect -5 34 -1 38
rect -92 -10 -88 -6
rect -5 -10 -1 -6
rect -92 -54 -88 -50
rect -5 -54 -1 -50
<< ntransistor >>
rect -92 0 -72 2
rect 0 0 4 2
rect -92 -18 -72 -16
rect 0 -18 4 -16
rect 0 -22 4 -20
<< ptransistor >>
rect -92 26 -72 28
rect 0 26 4 28
rect -92 -44 -72 -42
rect 0 -44 4 -42
rect 10 -44 14 -42
<< psubstratepcontact >>
rect -87 -11 -83 -5
rect 0 -11 4 -5
<< nsubstratencontact >>
rect -87 33 -82 38
rect 0 33 5 38
rect -87 -54 -82 -49
rect 0 -54 5 -49
<< labels >>
rlabel metal2 -43 -8 -43 -8 1 GND!
rlabel metal2 -41 36 -41 36 5 Vdd!
rlabel metal2 -43 -8 -43 -8 5 GND!
rlabel metal2 -41 -52 -41 -52 1 Vdd!
rlabel polysilicon -37 -32 -37 -32 1 net2
rlabel polysilicon -36 16 -36 16 1 net1
rlabel metal1 -101 -32 -101 -32 3 in2
rlabel metal1 -101 16 -101 16 3 in1
rlabel metal1 2 12 2 12 1 out1
rlabel metal1 2 -30 2 -30 1 out2
<< end >>
