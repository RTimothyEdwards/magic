magic
tech nmos
timestamp 478544012
<< polysilicon >>
rect -10 8 -8 10
rect -6 8 10 10
rect -10 1 -8 5
rect -6 1 -3 5
<< diffusion >>
rect -8 10 -6 12
rect -8 5 -6 8
rect -8 -1 -6 1
rect -8 -9 -6 -5
<< metal >>
rect 1 1 10 4
rect -6 -5 10 -2
<< poly-metal-contact >>
rect -3 1 1 5
<< diff-metal-contact >>
rect -10 -5 -6 -1
<< enhancement-fet >>
rect -8 8 -6 10
<< depletion-fet >>
rect -8 1 -6 5
<< end >>
