magic
tech scmos
timestamp 500618582
<< polysilicon >>
rect 1 8 7 11
rect 5 5 7 8
rect -9 -6 -6 1
rect 2 -5 6 0
<< end >>
