magic
tech scmos
timestamp 616443648
<< polysilicon >>
rect -3 104 -1 106
rect 38 104 40 106
rect -3 96 -1 101
rect -3 94 7 96
rect -9 88 -7 90
rect 9 88 11 94
rect 25 94 26 96
rect 38 96 40 101
rect 30 94 40 96
rect 25 88 27 94
rect 44 88 46 90
rect -3 81 -1 83
rect -9 79 -7 80
rect 38 81 40 83
rect 44 79 46 80
<< ndiffusion >>
rect -12 86 -9 88
rect -11 82 -9 86
rect -12 80 -9 82
rect -7 84 -1 88
rect 3 84 9 88
rect -7 80 -4 84
rect -1 83 9 84
rect 11 83 25 88
rect 27 84 34 88
rect 38 84 44 88
rect 27 83 38 84
rect 11 81 14 83
rect -1 79 14 81
rect 24 81 25 83
rect 24 79 38 81
rect 41 80 44 84
rect 46 80 49 88
rect -1 78 18 79
rect 23 78 38 79
<< pdiffusion >>
rect -8 108 1 112
rect 36 108 45 112
rect -8 104 -4 108
rect 41 104 45 108
rect -8 101 -3 104
rect -1 101 0 104
rect 37 101 38 104
rect 40 101 45 104
<< metal1 >>
rect -12 99 -9 112
rect -6 105 -3 112
rect -6 104 3 105
rect -6 102 0 104
rect -12 96 -5 99
rect -12 89 -11 92
rect -16 86 -11 89
rect -8 79 -5 96
rect 0 88 3 100
rect 8 99 11 112
rect 14 91 17 112
rect 7 88 17 91
rect 20 91 23 112
rect 26 99 29 112
rect 40 104 43 112
rect 37 101 43 104
rect 20 88 30 91
rect -6 74 -5 79
rect -8 72 -5 74
rect 7 72 10 88
rect 14 78 24 79
rect 18 77 23 78
rect 18 74 19 77
rect 27 72 30 88
rect 34 88 37 100
rect 46 98 49 112
rect 42 95 49 98
rect 42 79 45 95
rect 42 74 43 79
rect 42 72 45 74
<< metal2 >>
rect -16 93 55 97
rect -12 89 -11 93
rect -16 86 -11 89
rect -16 77 55 79
rect -16 74 19 77
rect 23 74 55 77
<< polycontact >>
rect 7 94 11 99
rect 26 94 30 99
rect -11 74 -6 79
rect 43 74 48 79
<< ndcontact >>
rect -16 82 -11 86
rect -1 84 3 88
rect 34 84 38 88
rect 14 79 24 83
<< pdcontact >>
rect 0 100 4 104
rect 33 100 37 104
<< m2contact >>
rect -16 89 -12 93
rect 19 73 23 77
<< ntransistor >>
rect -9 80 -7 88
rect 9 83 11 88
rect 25 83 27 88
rect -1 81 11 83
rect 25 81 38 83
rect 44 80 46 88
<< ptransistor >>
rect -3 101 -1 104
rect 38 101 40 104
<< psubstratepcontact >>
rect 13 74 18 78
<< nsubstratencontact >>
rect 1 108 5 112
rect 32 108 36 112
<< labels >>
rlabel metal1 -8 72 -5 72 1 accA0
rlabel metal1 7 72 10 72 1 accB0
rlabel metal1 27 72 30 72 1 accB1
rlabel metal1 42 72 45 72 1 accA1
rlabel metal2 55 74 55 79 7 GND!
rlabel metal2 55 93 55 97 7 busA0
<< end >>
